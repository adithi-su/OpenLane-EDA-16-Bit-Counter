magic
tech sky130A
magscale 1 2
timestamp 1647516069
<< obsli1 >>
rect 1104 2159 13800 14705
<< obsm1 >>
rect 14 2128 14890 14736
<< metal2 >>
rect 2594 16325 2650 17125
rect 5814 16325 5870 17125
rect 9034 16325 9090 17125
rect 12254 16325 12310 17125
rect 14830 16325 14886 17125
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 9034 0 9090 800
rect 12254 0 12310 800
<< obsm2 >>
rect 20 16269 2538 16425
rect 2706 16269 5758 16425
rect 5926 16269 8978 16425
rect 9146 16269 12198 16425
rect 12366 16269 14774 16425
rect 20 856 14884 16269
rect 130 31 2538 856
rect 2706 31 5758 856
rect 5926 31 8978 856
rect 9146 31 12198 856
rect 12366 31 14884 856
<< metal3 >>
rect 0 16328 800 16448
rect 14181 13608 14981 13728
rect 0 12928 800 13048
rect 14181 10208 14981 10328
rect 0 9528 800 9648
rect 14181 6808 14981 6928
rect 0 6128 800 6248
rect 14181 3408 14981 3528
rect 0 2728 800 2848
rect 14181 8 14981 128
<< obsm3 >>
rect 880 16248 14181 16421
rect 800 13808 14181 16248
rect 800 13528 14101 13808
rect 800 13128 14181 13528
rect 880 12848 14181 13128
rect 800 10408 14181 12848
rect 800 10128 14101 10408
rect 800 9728 14181 10128
rect 880 9448 14181 9728
rect 800 7008 14181 9448
rect 800 6728 14101 7008
rect 800 6328 14181 6728
rect 880 6048 14181 6328
rect 800 3608 14181 6048
rect 800 3328 14101 3608
rect 800 2928 14181 3328
rect 880 2648 14181 2928
rect 800 208 14181 2648
rect 800 35 14101 208
<< metal4 >>
rect 3060 2128 3380 14736
rect 5176 2128 5496 14736
rect 7292 2128 7612 14736
rect 9408 2128 9728 14736
rect 11524 2128 11844 14736
<< metal5 >>
rect 1104 12395 13800 12715
rect 1104 10309 13800 10629
rect 1104 8224 13800 8544
rect 1104 6139 13800 6459
rect 1104 4053 13800 4373
<< obsm5 >>
rect 1104 10949 13800 12075
rect 1104 8864 13800 9989
rect 1104 6779 13800 7904
<< labels >>
rlabel metal5 s 1104 6139 13800 6459 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 10309 13800 10629 6 VGND
port 1 nsew ground input
rlabel metal4 s 5176 2128 5496 14736 6 VGND
port 1 nsew ground input
rlabel metal4 s 9408 2128 9728 14736 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 4053 13800 4373 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 8224 13800 8544 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 12395 13800 12715 6 VPWR
port 2 nsew power input
rlabel metal4 s 3060 2128 3380 14736 6 VPWR
port 2 nsew power input
rlabel metal4 s 7292 2128 7612 14736 6 VPWR
port 2 nsew power input
rlabel metal4 s 11524 2128 11844 14736 6 VPWR
port 2 nsew power input
rlabel metal3 s 14181 3408 14981 3528 6 clock
port 3 nsew signal input
rlabel metal2 s 14830 16325 14886 17125 6 count[0]
port 4 nsew signal output
rlabel metal2 s 9034 16325 9090 17125 6 count[10]
port 5 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 count[11]
port 6 nsew signal output
rlabel metal3 s 14181 13608 14981 13728 6 count[12]
port 7 nsew signal output
rlabel metal3 s 14181 8 14981 128 6 count[13]
port 8 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 count[14]
port 9 nsew signal output
rlabel metal2 s 5814 16325 5870 17125 6 count[15]
port 10 nsew signal output
rlabel metal2 s 18 0 74 800 6 count[1]
port 11 nsew signal output
rlabel metal2 s 2594 16325 2650 17125 6 count[2]
port 12 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 count[3]
port 13 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 count[4]
port 14 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 count[5]
port 15 nsew signal output
rlabel metal3 s 14181 10208 14981 10328 6 count[6]
port 16 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 count[7]
port 17 nsew signal output
rlabel metal2 s 12254 16325 12310 17125 6 count[8]
port 18 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 count[9]
port 19 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 count_en
port 20 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 count_tc
port 21 nsew signal output
rlabel metal3 s 14181 6808 14981 6928 6 reset
port 22 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 14981 17125
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 455626
string GDS_FILE /openlane/designs/counter_16b/runs/RUN_2022.03.17_11.20.16/results/finishing/counter_16b.magic.gds
string GDS_START 159472
<< end >>

