magic
tech sky130A
magscale 1 2
timestamp 1647516074
<< checkpaint >>
rect -3932 -3932 18913 21057
<< viali >>
rect 1501 14569 1535 14603
rect 2789 14569 2823 14603
rect 6561 14569 6595 14603
rect 9229 14569 9263 14603
rect 12265 14569 12299 14603
rect 13001 14569 13035 14603
rect 1685 14365 1719 14399
rect 2973 14365 3007 14399
rect 6377 14365 6411 14399
rect 9413 14365 9447 14399
rect 12081 14365 12115 14399
rect 12817 14365 12851 14399
rect 12817 13889 12851 13923
rect 13001 13685 13035 13719
rect 1685 13277 1719 13311
rect 1501 13141 1535 13175
rect 6561 11645 6595 11679
rect 6929 11577 6963 11611
rect 7021 11509 7055 11543
rect 7297 11305 7331 11339
rect 4813 11169 4847 11203
rect 8125 11169 8159 11203
rect 8401 11169 8435 11203
rect 1409 11101 1443 11135
rect 4905 11101 4939 11135
rect 4997 11101 5031 11135
rect 5917 11101 5951 11135
rect 7941 11101 7975 11135
rect 8033 11101 8067 11135
rect 8217 11101 8251 11135
rect 6184 11033 6218 11067
rect 1593 10965 1627 10999
rect 4629 10965 4663 10999
rect 5089 10761 5123 10795
rect 5641 10761 5675 10795
rect 6745 10761 6779 10795
rect 6653 10693 6687 10727
rect 7649 10693 7683 10727
rect 7849 10693 7883 10727
rect 1777 10625 1811 10659
rect 2044 10625 2078 10659
rect 3709 10625 3743 10659
rect 3965 10625 3999 10659
rect 5825 10625 5859 10659
rect 6469 10625 6503 10659
rect 6837 10625 6871 10659
rect 8309 10625 8343 10659
rect 12817 10625 12851 10659
rect 7021 10557 7055 10591
rect 8585 10557 8619 10591
rect 9597 10557 9631 10591
rect 7481 10489 7515 10523
rect 9873 10489 9907 10523
rect 3157 10421 3191 10455
rect 7665 10421 7699 10455
rect 10057 10421 10091 10455
rect 13001 10421 13035 10455
rect 1961 10217 1995 10251
rect 2329 10217 2363 10251
rect 5917 10217 5951 10251
rect 6469 10217 6503 10251
rect 7113 10217 7147 10251
rect 10333 10217 10367 10251
rect 2881 10149 2915 10183
rect 4537 10081 4571 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 2145 10013 2179 10047
rect 2421 10013 2455 10047
rect 3065 10013 3099 10047
rect 3157 10013 3191 10047
rect 4793 10013 4827 10047
rect 6653 10013 6687 10047
rect 7757 10013 7791 10047
rect 8217 10013 8251 10047
rect 8953 10013 8987 10047
rect 2881 9945 2915 9979
rect 9220 9945 9254 9979
rect 7573 9877 7607 9911
rect 7665 9877 7699 9911
rect 8309 9877 8343 9911
rect 3801 9673 3835 9707
rect 4445 9673 4479 9707
rect 4261 9605 4295 9639
rect 2614 9537 2648 9571
rect 2881 9537 2915 9571
rect 3341 9537 3375 9571
rect 3617 9537 3651 9571
rect 4537 9537 4571 9571
rect 5457 9537 5491 9571
rect 5733 9537 5767 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 8677 9537 8711 9571
rect 8861 9537 8895 9571
rect 9588 9537 9622 9571
rect 5273 9469 5307 9503
rect 5549 9469 5583 9503
rect 5641 9469 5675 9503
rect 6377 9469 6411 9503
rect 6561 9469 6595 9503
rect 6653 9469 6687 9503
rect 7389 9469 7423 9503
rect 7665 9469 7699 9503
rect 9321 9469 9355 9503
rect 4261 9401 4295 9435
rect 1501 9333 1535 9367
rect 3433 9333 3467 9367
rect 8769 9333 8803 9367
rect 10701 9333 10735 9367
rect 2605 9129 2639 9163
rect 3985 9129 4019 9163
rect 4721 9129 4755 9163
rect 8217 9129 8251 9163
rect 9229 9129 9263 9163
rect 9689 9129 9723 9163
rect 6561 8993 6595 9027
rect 7941 8993 7975 9027
rect 1961 8925 1995 8959
rect 6285 8925 6319 8959
rect 7573 8925 7607 8959
rect 8033 8925 8067 8959
rect 8953 8925 8987 8959
rect 9045 8925 9079 8959
rect 9873 8925 9907 8959
rect 1685 8857 1719 8891
rect 1869 8857 1903 8891
rect 2421 8857 2455 8891
rect 2621 8857 2655 8891
rect 3801 8857 3835 8891
rect 4017 8857 4051 8891
rect 4813 8857 4847 8891
rect 9229 8857 9263 8891
rect 1783 8789 1817 8823
rect 2789 8789 2823 8823
rect 4169 8789 4203 8823
rect 7665 8789 7699 8823
rect 7849 8789 7883 8823
rect 2145 8585 2179 8619
rect 8309 8585 8343 8619
rect 2421 8517 2455 8551
rect 5549 8517 5583 8551
rect 2145 8449 2179 8483
rect 3341 8449 3375 8483
rect 4813 8449 4847 8483
rect 5457 8449 5491 8483
rect 5733 8449 5767 8483
rect 6653 8449 6687 8483
rect 7941 8449 7975 8483
rect 8125 8449 8159 8483
rect 8953 8449 8987 8483
rect 3617 8381 3651 8415
rect 4997 8381 5031 8415
rect 6377 8381 6411 8415
rect 7849 8381 7883 8415
rect 8033 8381 8067 8415
rect 2237 8313 2271 8347
rect 5733 8313 5767 8347
rect 8769 8313 8803 8347
rect 4629 8245 4663 8279
rect 5549 8041 5583 8075
rect 8217 8041 8251 8075
rect 2881 7905 2915 7939
rect 9321 7905 9355 7939
rect 3065 7837 3099 7871
rect 4169 7837 4203 7871
rect 6009 7837 6043 7871
rect 7849 7837 7883 7871
rect 4414 7769 4448 7803
rect 6254 7769 6288 7803
rect 9505 7769 9539 7803
rect 3249 7701 3283 7735
rect 7389 7701 7423 7735
rect 8217 7701 8251 7735
rect 8401 7701 8435 7735
rect 3893 7497 3927 7531
rect 4537 7497 4571 7531
rect 5825 7497 5859 7531
rect 8401 7497 8435 7531
rect 3617 7429 3651 7463
rect 4353 7429 4387 7463
rect 9597 7429 9631 7463
rect 2053 7361 2087 7395
rect 2881 7361 2915 7395
rect 3065 7361 3099 7395
rect 3801 7361 3835 7395
rect 3893 7361 3927 7395
rect 4629 7361 4663 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 5365 7361 5399 7395
rect 5641 7361 5675 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 7941 7361 7975 7395
rect 8585 7361 8619 7395
rect 8677 7361 8711 7395
rect 8769 7361 8803 7395
rect 9413 7361 9447 7395
rect 9689 7361 9723 7395
rect 12817 7361 12851 7395
rect 1961 7293 1995 7327
rect 2145 7293 2179 7327
rect 3157 7293 3191 7327
rect 6469 7293 6503 7327
rect 7665 7293 7699 7327
rect 8861 7293 8895 7327
rect 13093 7293 13127 7327
rect 1777 7157 1811 7191
rect 2697 7157 2731 7191
rect 5457 7157 5491 7191
rect 9413 7157 9447 7191
rect 4997 6953 5031 6987
rect 7113 6953 7147 6987
rect 8953 6953 8987 6987
rect 3801 6817 3835 6851
rect 4077 6817 4111 6851
rect 4261 6817 4295 6851
rect 8033 6817 8067 6851
rect 8125 6817 8159 6851
rect 1501 6749 1535 6783
rect 1768 6749 1802 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 6377 6749 6411 6783
rect 6469 6749 6503 6783
rect 7941 6749 7975 6783
rect 8217 6749 8251 6783
rect 10333 6749 10367 6783
rect 4965 6681 4999 6715
rect 5181 6681 5215 6715
rect 6193 6681 6227 6715
rect 6929 6681 6963 6715
rect 7145 6681 7179 6715
rect 10066 6681 10100 6715
rect 2881 6613 2915 6647
rect 4813 6613 4847 6647
rect 6291 6613 6325 6647
rect 7297 6613 7331 6647
rect 7757 6613 7791 6647
rect 1768 6341 1802 6375
rect 1501 6273 1535 6307
rect 4537 6273 4571 6307
rect 4997 6273 5031 6307
rect 5089 6273 5123 6307
rect 5273 6273 5307 6307
rect 6653 6273 6687 6307
rect 8421 6273 8455 6307
rect 9413 6273 9447 6307
rect 4261 6205 4295 6239
rect 6377 6205 6411 6239
rect 8677 6205 8711 6239
rect 9137 6205 9171 6239
rect 2881 6137 2915 6171
rect 5273 6069 5307 6103
rect 6469 6069 6503 6103
rect 6837 6069 6871 6103
rect 7297 6069 7331 6103
rect 1501 5865 1535 5899
rect 2329 5865 2363 5899
rect 8953 5865 8987 5899
rect 3801 5797 3835 5831
rect 4997 5729 5031 5763
rect 5089 5729 5123 5763
rect 5273 5729 5307 5763
rect 6929 5729 6963 5763
rect 1685 5661 1719 5695
rect 2145 5661 2179 5695
rect 2329 5661 2363 5695
rect 2789 5661 2823 5695
rect 3065 5661 3099 5695
rect 3985 5661 4019 5695
rect 5181 5661 5215 5695
rect 7185 5661 7219 5695
rect 9137 5661 9171 5695
rect 4169 5593 4203 5627
rect 4353 5593 4387 5627
rect 2881 5525 2915 5559
rect 3249 5525 3283 5559
rect 4077 5525 4111 5559
rect 4813 5525 4847 5559
rect 8309 5525 8343 5559
rect 8033 5321 8067 5355
rect 3065 5185 3099 5219
rect 4353 5185 4387 5219
rect 4620 5185 4654 5219
rect 7941 5185 7975 5219
rect 8125 5185 8159 5219
rect 3341 5117 3375 5151
rect 5733 5049 5767 5083
rect 4905 4777 4939 4811
rect 3985 4573 4019 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 4905 4573 4939 4607
rect 5089 4573 5123 4607
rect 3801 4437 3835 4471
rect 3648 4165 3682 4199
rect 3893 4097 3927 4131
rect 2513 3893 2547 3927
rect 12817 3553 12851 3587
rect 13093 3485 13127 3519
rect 1685 3009 1719 3043
rect 1501 2805 1535 2839
rect 13001 2533 13035 2567
rect 1685 2397 1719 2431
rect 2973 2397 3007 2431
rect 6653 2397 6687 2431
rect 9137 2397 9171 2431
rect 12081 2397 12115 2431
rect 12817 2397 12851 2431
rect 1501 2261 1535 2295
rect 2789 2261 2823 2295
rect 6469 2261 6503 2295
rect 9321 2261 9355 2295
rect 12265 2261 12299 2295
<< metal1 >>
rect 1104 14714 13800 14736
rect 1104 14662 3066 14714
rect 3118 14662 3130 14714
rect 3182 14662 3194 14714
rect 3246 14662 3258 14714
rect 3310 14662 3322 14714
rect 3374 14662 7298 14714
rect 7350 14662 7362 14714
rect 7414 14662 7426 14714
rect 7478 14662 7490 14714
rect 7542 14662 7554 14714
rect 7606 14662 11530 14714
rect 11582 14662 11594 14714
rect 11646 14662 11658 14714
rect 11710 14662 11722 14714
rect 11774 14662 11786 14714
rect 11838 14662 13800 14714
rect 1104 14640 13800 14662
rect 1486 14600 1492 14612
rect 1447 14572 1492 14600
rect 1486 14560 1492 14572
rect 1544 14560 1550 14612
rect 2774 14600 2780 14612
rect 2735 14572 2780 14600
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 6549 14603 6607 14609
rect 6549 14600 6561 14603
rect 5868 14572 6561 14600
rect 5868 14560 5874 14572
rect 6549 14569 6561 14572
rect 6595 14569 6607 14603
rect 6549 14563 6607 14569
rect 9030 14560 9036 14612
rect 9088 14600 9094 14612
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 9088 14572 9229 14600
rect 9088 14560 9094 14572
rect 9217 14569 9229 14572
rect 9263 14569 9275 14603
rect 12250 14600 12256 14612
rect 12211 14572 12256 14600
rect 9217 14563 9275 14569
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 12989 14603 13047 14609
rect 12989 14569 13001 14603
rect 13035 14600 13047 14603
rect 14826 14600 14832 14612
rect 13035 14572 14832 14600
rect 13035 14569 13047 14572
rect 12989 14563 13047 14569
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 4154 14396 4160 14408
rect 3007 14368 4160 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 1688 14328 1716 14359
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 5902 14356 5908 14408
rect 5960 14396 5966 14408
rect 6365 14399 6423 14405
rect 6365 14396 6377 14399
rect 5960 14368 6377 14396
rect 5960 14356 5966 14368
rect 6365 14365 6377 14368
rect 6411 14365 6423 14399
rect 6365 14359 6423 14365
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9364 14368 9413 14396
rect 9364 14356 9370 14368
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 12066 14396 12072 14408
rect 12027 14368 12072 14396
rect 9401 14359 9459 14365
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 12492 14368 12817 14396
rect 12492 14356 12498 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 4798 14328 4804 14340
rect 1688 14300 4804 14328
rect 4798 14288 4804 14300
rect 4856 14288 4862 14340
rect 1104 14170 13800 14192
rect 1104 14118 5182 14170
rect 5234 14118 5246 14170
rect 5298 14118 5310 14170
rect 5362 14118 5374 14170
rect 5426 14118 5438 14170
rect 5490 14118 9414 14170
rect 9466 14118 9478 14170
rect 9530 14118 9542 14170
rect 9594 14118 9606 14170
rect 9658 14118 9670 14170
rect 9722 14118 13800 14170
rect 1104 14096 13800 14118
rect 10318 13880 10324 13932
rect 10376 13920 10382 13932
rect 12805 13923 12863 13929
rect 12805 13920 12817 13923
rect 10376 13892 12817 13920
rect 10376 13880 10382 13892
rect 12805 13889 12817 13892
rect 12851 13889 12863 13923
rect 12805 13883 12863 13889
rect 12986 13716 12992 13728
rect 12947 13688 12992 13716
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 1104 13626 13800 13648
rect 1104 13574 3066 13626
rect 3118 13574 3130 13626
rect 3182 13574 3194 13626
rect 3246 13574 3258 13626
rect 3310 13574 3322 13626
rect 3374 13574 7298 13626
rect 7350 13574 7362 13626
rect 7414 13574 7426 13626
rect 7478 13574 7490 13626
rect 7542 13574 7554 13626
rect 7606 13574 11530 13626
rect 11582 13574 11594 13626
rect 11646 13574 11658 13626
rect 11710 13574 11722 13626
rect 11774 13574 11786 13626
rect 11838 13574 13800 13626
rect 1104 13552 13800 13574
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 7190 13308 7196 13320
rect 1719 13280 7196 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 1104 13082 13800 13104
rect 1104 13030 5182 13082
rect 5234 13030 5246 13082
rect 5298 13030 5310 13082
rect 5362 13030 5374 13082
rect 5426 13030 5438 13082
rect 5490 13030 9414 13082
rect 9466 13030 9478 13082
rect 9530 13030 9542 13082
rect 9594 13030 9606 13082
rect 9658 13030 9670 13082
rect 9722 13030 13800 13082
rect 1104 13008 13800 13030
rect 1104 12538 13800 12560
rect 1104 12486 3066 12538
rect 3118 12486 3130 12538
rect 3182 12486 3194 12538
rect 3246 12486 3258 12538
rect 3310 12486 3322 12538
rect 3374 12486 7298 12538
rect 7350 12486 7362 12538
rect 7414 12486 7426 12538
rect 7478 12486 7490 12538
rect 7542 12486 7554 12538
rect 7606 12486 11530 12538
rect 11582 12486 11594 12538
rect 11646 12486 11658 12538
rect 11710 12486 11722 12538
rect 11774 12486 11786 12538
rect 11838 12486 13800 12538
rect 1104 12464 13800 12486
rect 1104 11994 13800 12016
rect 1104 11942 5182 11994
rect 5234 11942 5246 11994
rect 5298 11942 5310 11994
rect 5362 11942 5374 11994
rect 5426 11942 5438 11994
rect 5490 11942 9414 11994
rect 9466 11942 9478 11994
rect 9530 11942 9542 11994
rect 9594 11942 9606 11994
rect 9658 11942 9670 11994
rect 9722 11942 13800 11994
rect 1104 11920 13800 11942
rect 6362 11636 6368 11688
rect 6420 11676 6426 11688
rect 6549 11679 6607 11685
rect 6549 11676 6561 11679
rect 6420 11648 6561 11676
rect 6420 11636 6426 11648
rect 6549 11645 6561 11648
rect 6595 11645 6607 11679
rect 6549 11639 6607 11645
rect 6914 11608 6920 11620
rect 6875 11580 6920 11608
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7006 11540 7012 11552
rect 6967 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 1104 11450 13800 11472
rect 1104 11398 3066 11450
rect 3118 11398 3130 11450
rect 3182 11398 3194 11450
rect 3246 11398 3258 11450
rect 3310 11398 3322 11450
rect 3374 11398 7298 11450
rect 7350 11398 7362 11450
rect 7414 11398 7426 11450
rect 7478 11398 7490 11450
rect 7542 11398 7554 11450
rect 7606 11398 11530 11450
rect 11582 11398 11594 11450
rect 11646 11398 11658 11450
rect 11710 11398 11722 11450
rect 11774 11398 11786 11450
rect 11838 11398 13800 11450
rect 1104 11376 13800 11398
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 7248 11308 7297 11336
rect 7248 11296 7254 11308
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 7285 11299 7343 11305
rect 4798 11200 4804 11212
rect 4759 11172 4804 11200
rect 4798 11160 4804 11172
rect 4856 11200 4862 11212
rect 5626 11200 5632 11212
rect 4856 11172 5632 11200
rect 4856 11160 4862 11172
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 8110 11200 8116 11212
rect 8071 11172 8116 11200
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 9858 11200 9864 11212
rect 8435 11172 9864 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 9858 11160 9864 11172
rect 9916 11160 9922 11212
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 4890 11132 4896 11144
rect 4851 11104 4896 11132
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 5905 11135 5963 11141
rect 5040 11104 5085 11132
rect 5040 11092 5046 11104
rect 5905 11101 5917 11135
rect 5951 11101 5963 11135
rect 7926 11132 7932 11144
rect 7887 11104 7932 11132
rect 5905 11095 5963 11101
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5920 11064 5948 11095
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 5132 11036 5948 11064
rect 6172 11067 6230 11073
rect 5132 11024 5138 11036
rect 6172 11033 6184 11067
rect 6218 11064 6230 11067
rect 6454 11064 6460 11076
rect 6218 11036 6460 11064
rect 6218 11033 6230 11036
rect 6172 11027 6230 11033
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 8036 11064 8064 11095
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8260 11104 8305 11132
rect 8260 11092 8266 11104
rect 8036 11036 8248 11064
rect 8220 11008 8248 11036
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10996 1639 10999
rect 2406 10996 2412 11008
rect 1627 10968 2412 10996
rect 1627 10965 1639 10968
rect 1581 10959 1639 10965
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 4614 10996 4620 11008
rect 4575 10968 4620 10996
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 8202 10956 8208 11008
rect 8260 10956 8266 11008
rect 1104 10906 13800 10928
rect 1104 10854 5182 10906
rect 5234 10854 5246 10906
rect 5298 10854 5310 10906
rect 5362 10854 5374 10906
rect 5426 10854 5438 10906
rect 5490 10854 9414 10906
rect 9466 10854 9478 10906
rect 9530 10854 9542 10906
rect 9594 10854 9606 10906
rect 9658 10854 9670 10906
rect 9722 10854 13800 10906
rect 1104 10832 13800 10854
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 5077 10795 5135 10801
rect 5077 10792 5089 10795
rect 4212 10764 5089 10792
rect 4212 10752 4218 10764
rect 5077 10761 5089 10764
rect 5123 10761 5135 10795
rect 5626 10792 5632 10804
rect 5587 10764 5632 10792
rect 5077 10755 5135 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 6733 10795 6791 10801
rect 6733 10761 6745 10795
rect 6779 10792 6791 10795
rect 7098 10792 7104 10804
rect 6779 10764 7104 10792
rect 6779 10761 6791 10764
rect 6733 10755 6791 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7248 10764 7880 10792
rect 7248 10752 7254 10764
rect 2866 10724 2872 10736
rect 1780 10696 2872 10724
rect 1780 10665 1808 10696
rect 2866 10684 2872 10696
rect 2924 10724 2930 10736
rect 2924 10696 5120 10724
rect 2924 10684 2930 10696
rect 2038 10665 2044 10668
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 2032 10619 2044 10665
rect 2096 10656 2102 10668
rect 3712 10665 3740 10696
rect 5092 10668 5120 10696
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 7852 10733 7880 10764
rect 6641 10727 6699 10733
rect 6641 10724 6653 10727
rect 6604 10696 6653 10724
rect 6604 10684 6610 10696
rect 6641 10693 6653 10696
rect 6687 10724 6699 10727
rect 7637 10727 7695 10733
rect 6687 10696 7512 10724
rect 6687 10693 6699 10696
rect 6641 10687 6699 10693
rect 3697 10659 3755 10665
rect 2096 10628 2132 10656
rect 2038 10616 2044 10619
rect 2096 10616 2102 10628
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3953 10659 4011 10665
rect 3953 10656 3965 10659
rect 3844 10628 3965 10656
rect 3844 10616 3850 10628
rect 3953 10625 3965 10628
rect 3999 10625 4011 10659
rect 3953 10619 4011 10625
rect 5074 10616 5080 10668
rect 5132 10616 5138 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6457 10659 6515 10665
rect 6457 10656 6469 10659
rect 5859 10628 6469 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6457 10625 6469 10628
rect 6503 10625 6515 10659
rect 6457 10619 6515 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 7374 10656 7380 10668
rect 6871 10628 7380 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 5960 10560 7021 10588
rect 5960 10548 5966 10560
rect 7009 10557 7021 10560
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7484 10529 7512 10696
rect 7637 10693 7649 10727
rect 7683 10724 7695 10727
rect 7837 10727 7895 10733
rect 7683 10696 7788 10724
rect 7683 10693 7695 10696
rect 7637 10687 7695 10693
rect 7760 10656 7788 10696
rect 7837 10693 7849 10727
rect 7883 10693 7895 10727
rect 7837 10687 7895 10693
rect 8297 10659 8355 10665
rect 8297 10656 8309 10659
rect 7760 10628 8309 10656
rect 8297 10625 8309 10628
rect 8343 10656 8355 10659
rect 10318 10656 10324 10668
rect 8343 10628 10324 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12676 10628 12817 10656
rect 12676 10616 12682 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8260 10560 8585 10588
rect 8260 10548 8266 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 8812 10560 9597 10588
rect 8812 10548 8818 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 12434 10588 12440 10600
rect 9585 10551 9643 10557
rect 9692 10560 12440 10588
rect 7469 10523 7527 10529
rect 5000 10492 5396 10520
rect 3145 10455 3203 10461
rect 3145 10421 3157 10455
rect 3191 10452 3203 10455
rect 3418 10452 3424 10464
rect 3191 10424 3424 10452
rect 3191 10421 3203 10424
rect 3145 10415 3203 10421
rect 3418 10412 3424 10424
rect 3476 10452 3482 10464
rect 5000 10452 5028 10492
rect 3476 10424 5028 10452
rect 5368 10452 5396 10492
rect 7469 10489 7481 10523
rect 7515 10489 7527 10523
rect 9692 10520 9720 10560
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 9858 10520 9864 10532
rect 7469 10483 7527 10489
rect 7576 10492 9720 10520
rect 9819 10492 9864 10520
rect 7576 10452 7604 10492
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 5368 10424 7604 10452
rect 7653 10455 7711 10461
rect 3476 10412 3482 10424
rect 7653 10421 7665 10455
rect 7699 10452 7711 10455
rect 7926 10452 7932 10464
rect 7699 10424 7932 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 1104 10362 13800 10384
rect 1104 10310 3066 10362
rect 3118 10310 3130 10362
rect 3182 10310 3194 10362
rect 3246 10310 3258 10362
rect 3310 10310 3322 10362
rect 3374 10310 7298 10362
rect 7350 10310 7362 10362
rect 7414 10310 7426 10362
rect 7478 10310 7490 10362
rect 7542 10310 7554 10362
rect 7606 10310 11530 10362
rect 11582 10310 11594 10362
rect 11646 10310 11658 10362
rect 11710 10310 11722 10362
rect 11774 10310 11786 10362
rect 11838 10310 13800 10362
rect 1104 10288 13800 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2038 10248 2044 10260
rect 1995 10220 2044 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2590 10248 2596 10260
rect 2363 10220 2596 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2590 10208 2596 10220
rect 2648 10248 2654 10260
rect 5166 10248 5172 10260
rect 2648 10220 3188 10248
rect 2648 10208 2654 10220
rect 2869 10183 2927 10189
rect 2869 10180 2881 10183
rect 2746 10152 2881 10180
rect 2746 10112 2774 10152
rect 2869 10149 2881 10152
rect 2915 10149 2927 10183
rect 2869 10143 2927 10149
rect 2148 10084 2774 10112
rect 2148 10053 2176 10084
rect 2133 10047 2191 10053
rect 2133 10013 2145 10047
rect 2179 10013 2191 10047
rect 2133 10007 2191 10013
rect 2406 10004 2412 10056
rect 2464 10044 2470 10056
rect 3160 10053 3188 10220
rect 4540 10220 5172 10248
rect 4540 10121 4568 10220
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5902 10248 5908 10260
rect 5863 10220 5908 10248
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 6454 10248 6460 10260
rect 6415 10220 6460 10248
rect 6454 10208 6460 10220
rect 6512 10208 6518 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 6972 10220 7113 10248
rect 6972 10208 6978 10220
rect 7101 10217 7113 10220
rect 7147 10217 7159 10251
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 7101 10211 7159 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 7248 10084 7297 10112
rect 7248 10072 7254 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7926 10112 7932 10124
rect 7423 10084 7932 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 2464 10016 3065 10044
rect 2464 10004 2470 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3418 10044 3424 10056
rect 3191 10016 3424 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 4781 10047 4839 10053
rect 4781 10044 4793 10047
rect 4672 10016 4793 10044
rect 4672 10004 4678 10016
rect 4781 10013 4793 10016
rect 4827 10013 4839 10047
rect 4781 10007 4839 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 7006 10044 7012 10056
rect 6687 10016 7012 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7708 10016 7757 10044
rect 7708 10004 7714 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 8202 10044 8208 10056
rect 8163 10016 8208 10044
rect 7745 10007 7803 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10044 8999 10047
rect 9030 10044 9036 10056
rect 8987 10016 9036 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 2869 9979 2927 9985
rect 2869 9976 2881 9979
rect 2740 9948 2881 9976
rect 2740 9936 2746 9948
rect 2869 9945 2881 9948
rect 2915 9976 2927 9979
rect 4890 9976 4896 9988
rect 2915 9948 4896 9976
rect 2915 9945 2927 9948
rect 2869 9939 2927 9945
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 7834 9976 7840 9988
rect 7576 9948 7840 9976
rect 7576 9917 7604 9948
rect 7834 9936 7840 9948
rect 7892 9976 7898 9988
rect 8220 9976 8248 10004
rect 9214 9985 9220 9988
rect 9208 9976 9220 9985
rect 7892 9948 8248 9976
rect 9175 9948 9220 9976
rect 7892 9936 7898 9948
rect 9208 9939 9220 9948
rect 9214 9936 9220 9939
rect 9272 9936 9278 9988
rect 7561 9911 7619 9917
rect 7561 9877 7573 9911
rect 7607 9877 7619 9911
rect 7561 9871 7619 9877
rect 7653 9911 7711 9917
rect 7653 9877 7665 9911
rect 7699 9908 7711 9911
rect 7742 9908 7748 9920
rect 7699 9880 7748 9908
rect 7699 9877 7711 9880
rect 7653 9871 7711 9877
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 9030 9908 9036 9920
rect 8343 9880 9036 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 1104 9818 13800 9840
rect 1104 9766 5182 9818
rect 5234 9766 5246 9818
rect 5298 9766 5310 9818
rect 5362 9766 5374 9818
rect 5426 9766 5438 9818
rect 5490 9766 9414 9818
rect 9466 9766 9478 9818
rect 9530 9766 9542 9818
rect 9594 9766 9606 9818
rect 9658 9766 9670 9818
rect 9722 9766 13800 9818
rect 1104 9744 13800 9766
rect 3786 9704 3792 9716
rect 3747 9676 3792 9704
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 4212 9676 4445 9704
rect 4212 9664 4218 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 4433 9667 4491 9673
rect 4172 9636 4200 9664
rect 3344 9608 4200 9636
rect 4249 9639 4307 9645
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2602 9571 2660 9577
rect 2602 9568 2614 9571
rect 2188 9540 2614 9568
rect 2188 9528 2194 9540
rect 2602 9537 2614 9540
rect 2648 9537 2660 9571
rect 2866 9568 2872 9580
rect 2827 9540 2872 9568
rect 2602 9531 2660 9537
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 3344 9577 3372 9608
rect 4249 9605 4261 9639
rect 4295 9636 4307 9639
rect 6546 9636 6552 9648
rect 4295 9608 5396 9636
rect 4295 9605 4307 9608
rect 4249 9599 4307 9605
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 3620 9500 3648 9531
rect 4540 9500 4568 9531
rect 3620 9472 4292 9500
rect 4264 9441 4292 9472
rect 4448 9472 4568 9500
rect 4249 9435 4307 9441
rect 4249 9401 4261 9435
rect 4295 9401 4307 9435
rect 4249 9395 4307 9401
rect 1489 9367 1547 9373
rect 1489 9333 1501 9367
rect 1535 9364 1547 9367
rect 1670 9364 1676 9376
rect 1535 9336 1676 9364
rect 1535 9333 1547 9336
rect 1489 9327 1547 9333
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 3421 9367 3479 9373
rect 3421 9333 3433 9367
rect 3467 9364 3479 9367
rect 3786 9364 3792 9376
rect 3467 9336 3792 9364
rect 3467 9333 3479 9336
rect 3421 9327 3479 9333
rect 3786 9324 3792 9336
rect 3844 9364 3850 9376
rect 4448 9364 4476 9472
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5040 9472 5273 9500
rect 5040 9460 5046 9472
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5261 9463 5319 9469
rect 3844 9336 4476 9364
rect 5368 9364 5396 9608
rect 5460 9608 6552 9636
rect 5460 9577 5488 9608
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 6914 9636 6920 9648
rect 6748 9608 6920 9636
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9568 5779 9571
rect 5902 9568 5908 9580
rect 5767 9540 5908 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 6748 9577 6776 9608
rect 6914 9596 6920 9608
rect 6972 9636 6978 9648
rect 8018 9636 8024 9648
rect 6972 9608 8024 9636
rect 6972 9596 6978 9608
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8168 9608 8708 9636
rect 8168 9596 8174 9608
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 6196 9540 6745 9568
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 6196 9500 6224 9540
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 8386 9568 8392 9580
rect 6871 9540 8392 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8680 9577 8708 9608
rect 9582 9577 9588 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 9576 9531 9588 9577
rect 9640 9568 9646 9580
rect 9640 9540 9676 9568
rect 6362 9500 6368 9512
rect 5675 9472 6224 9500
rect 6323 9472 6368 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 5552 9432 5580 9463
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 6546 9500 6552 9512
rect 6507 9472 6552 9500
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9469 6699 9503
rect 6641 9463 6699 9469
rect 6656 9432 6684 9463
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 7156 9472 7389 9500
rect 7156 9460 7162 9472
rect 7377 9469 7389 9472
rect 7423 9500 7435 9503
rect 7558 9500 7564 9512
rect 7423 9472 7564 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 8110 9500 8116 9512
rect 7699 9472 8116 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 7668 9432 7696 9463
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 8864 9500 8892 9531
rect 9582 9528 9588 9531
rect 9640 9528 9646 9540
rect 8260 9472 8892 9500
rect 8260 9460 8266 9472
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 9180 9472 9321 9500
rect 9180 9460 9186 9472
rect 9309 9469 9321 9472
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 5552 9404 7696 9432
rect 7926 9392 7932 9444
rect 7984 9432 7990 9444
rect 7984 9404 9076 9432
rect 7984 9392 7990 9404
rect 6362 9364 6368 9376
rect 5368 9336 6368 9364
rect 3844 9324 3850 9336
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8202 9364 8208 9376
rect 8076 9336 8208 9364
rect 8076 9324 8082 9336
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8757 9367 8815 9373
rect 8757 9333 8769 9367
rect 8803 9364 8815 9367
rect 8938 9364 8944 9376
rect 8803 9336 8944 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9048 9364 9076 9404
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 9048 9336 10701 9364
rect 10689 9333 10701 9336
rect 10735 9364 10747 9367
rect 12434 9364 12440 9376
rect 10735 9336 12440 9364
rect 10735 9333 10747 9336
rect 10689 9327 10747 9333
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 1104 9274 13800 9296
rect 1104 9222 3066 9274
rect 3118 9222 3130 9274
rect 3182 9222 3194 9274
rect 3246 9222 3258 9274
rect 3310 9222 3322 9274
rect 3374 9222 7298 9274
rect 7350 9222 7362 9274
rect 7414 9222 7426 9274
rect 7478 9222 7490 9274
rect 7542 9222 7554 9274
rect 7606 9222 11530 9274
rect 11582 9222 11594 9274
rect 11646 9222 11658 9274
rect 11710 9222 11722 9274
rect 11774 9222 11786 9274
rect 11838 9222 13800 9274
rect 1104 9200 13800 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 2593 9163 2651 9169
rect 2593 9160 2605 9163
rect 1728 9132 2605 9160
rect 1728 9120 1734 9132
rect 2593 9129 2605 9132
rect 2639 9129 2651 9163
rect 2593 9123 2651 9129
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 4614 9160 4620 9172
rect 4019 9132 4620 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9160 4767 9163
rect 4890 9160 4896 9172
rect 4755 9132 4896 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 8205 9163 8263 9169
rect 8205 9129 8217 9163
rect 8251 9160 8263 9163
rect 8754 9160 8760 9172
rect 8251 9132 8760 9160
rect 8251 9129 8263 9132
rect 8205 9123 8263 9129
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 9214 9160 9220 9172
rect 9175 9132 9220 9160
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9640 9132 9689 9160
rect 9640 9120 9646 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 9024 6607 9027
rect 6914 9024 6920 9036
rect 6595 8996 6920 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7926 9024 7932 9036
rect 7887 8996 7932 9024
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 6270 8956 6276 8968
rect 1995 8928 2636 8956
rect 6231 8928 6276 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2608 8900 2636 8928
rect 6270 8916 6276 8928
rect 6328 8916 6334 8968
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8956 7619 8959
rect 7650 8956 7656 8968
rect 7607 8928 7656 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8956 8079 8959
rect 8386 8956 8392 8968
rect 8067 8928 8392 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8938 8956 8944 8968
rect 8899 8928 8944 8956
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9861 8959 9919 8965
rect 9088 8928 9133 8956
rect 9088 8916 9094 8928
rect 9861 8925 9873 8959
rect 9907 8956 9919 8959
rect 10042 8956 10048 8968
rect 9907 8928 10048 8956
rect 9907 8925 9919 8928
rect 9861 8919 9919 8925
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 1670 8888 1676 8900
rect 1631 8860 1676 8888
rect 1670 8848 1676 8860
rect 1728 8848 1734 8900
rect 1857 8891 1915 8897
rect 1857 8857 1869 8891
rect 1903 8888 1915 8891
rect 2406 8888 2412 8900
rect 1903 8860 2412 8888
rect 1903 8857 1915 8860
rect 1857 8851 1915 8857
rect 2406 8848 2412 8860
rect 2464 8848 2470 8900
rect 2590 8848 2596 8900
rect 2648 8897 2654 8900
rect 2648 8891 2667 8897
rect 2655 8857 2667 8891
rect 3786 8888 3792 8900
rect 3747 8860 3792 8888
rect 2648 8851 2667 8857
rect 2648 8848 2654 8851
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 4005 8891 4063 8897
rect 4005 8857 4017 8891
rect 4051 8888 4063 8891
rect 4522 8888 4528 8900
rect 4051 8860 4528 8888
rect 4051 8857 4063 8860
rect 4005 8851 4063 8857
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 4798 8888 4804 8900
rect 4759 8860 4804 8888
rect 4798 8848 4804 8860
rect 4856 8848 4862 8900
rect 7742 8888 7748 8900
rect 7668 8860 7748 8888
rect 1762 8820 1768 8832
rect 1820 8829 1826 8832
rect 1729 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8783 1829 8829
rect 2777 8823 2835 8829
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 2866 8820 2872 8832
rect 2823 8792 2872 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 1820 8780 1826 8783
rect 2866 8780 2872 8792
rect 2924 8820 2930 8832
rect 3326 8820 3332 8832
rect 2924 8792 3332 8820
rect 2924 8780 2930 8792
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4246 8820 4252 8832
rect 4203 8792 4252 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 7668 8829 7696 8860
rect 7742 8848 7748 8860
rect 7800 8848 7806 8900
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 9217 8891 9275 8897
rect 9217 8888 9229 8891
rect 8352 8860 9229 8888
rect 8352 8848 8358 8860
rect 9217 8857 9229 8860
rect 9263 8857 9275 8891
rect 9217 8851 9275 8857
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8789 7711 8823
rect 7834 8820 7840 8832
rect 7795 8792 7840 8820
rect 7653 8783 7711 8789
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 1104 8730 13800 8752
rect 1104 8678 5182 8730
rect 5234 8678 5246 8730
rect 5298 8678 5310 8730
rect 5362 8678 5374 8730
rect 5426 8678 5438 8730
rect 5490 8678 9414 8730
rect 9466 8678 9478 8730
rect 9530 8678 9542 8730
rect 9594 8678 9606 8730
rect 9658 8678 9670 8730
rect 9722 8678 13800 8730
rect 1104 8656 13800 8678
rect 2130 8616 2136 8628
rect 2091 8588 2136 8616
rect 2130 8576 2136 8588
rect 2188 8576 2194 8628
rect 8294 8616 8300 8628
rect 8255 8588 8300 8616
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 2038 8508 2044 8560
rect 2096 8548 2102 8560
rect 2409 8551 2467 8557
rect 2409 8548 2421 8551
rect 2096 8520 2421 8548
rect 2096 8508 2102 8520
rect 2409 8517 2421 8520
rect 2455 8548 2467 8551
rect 2682 8548 2688 8560
rect 2455 8520 2688 8548
rect 2455 8517 2467 8520
rect 2409 8511 2467 8517
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 5537 8551 5595 8557
rect 5537 8548 5549 8551
rect 4816 8520 5549 8548
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 2133 8483 2191 8489
rect 2133 8480 2145 8483
rect 1820 8452 2145 8480
rect 1820 8440 1826 8452
rect 2133 8449 2145 8452
rect 2179 8449 2191 8483
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 2133 8443 2191 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4816 8489 4844 8520
rect 5537 8517 5549 8520
rect 5583 8517 5595 8551
rect 5537 8511 5595 8517
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 7892 8520 7972 8548
rect 7892 8508 7898 8520
rect 4801 8483 4859 8489
rect 4801 8480 4813 8483
rect 4212 8452 4813 8480
rect 4212 8440 4218 8452
rect 4801 8449 4813 8452
rect 4847 8449 4859 8483
rect 5445 8483 5503 8489
rect 5445 8480 5457 8483
rect 4801 8443 4859 8449
rect 4908 8452 5457 8480
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 3786 8412 3792 8424
rect 3651 8384 3792 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 2225 8347 2283 8353
rect 2225 8313 2237 8347
rect 2271 8344 2283 8347
rect 3620 8344 3648 8375
rect 3786 8372 3792 8384
rect 3844 8412 3850 8424
rect 4908 8412 4936 8452
rect 5445 8449 5457 8452
rect 5491 8449 5503 8483
rect 5718 8480 5724 8492
rect 5679 8452 5724 8480
rect 5445 8443 5503 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 7742 8480 7748 8492
rect 6687 8452 7748 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 7944 8489 7972 8520
rect 7929 8483 7987 8489
rect 7929 8449 7941 8483
rect 7975 8449 7987 8483
rect 8110 8480 8116 8492
rect 8071 8452 8116 8480
rect 7929 8443 7987 8449
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 8444 8452 8953 8480
rect 8444 8440 8450 8452
rect 8941 8449 8953 8452
rect 8987 8480 8999 8483
rect 9490 8480 9496 8492
rect 8987 8452 9496 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 3844 8384 4936 8412
rect 4985 8415 5043 8421
rect 3844 8372 3850 8384
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 5736 8412 5764 8440
rect 5031 8384 5764 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 6270 8372 6276 8424
rect 6328 8412 6334 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6328 8384 6377 8412
rect 6328 8372 6334 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 7837 8415 7895 8421
rect 7837 8381 7849 8415
rect 7883 8381 7895 8415
rect 8018 8412 8024 8424
rect 7979 8384 8024 8412
rect 7837 8375 7895 8381
rect 2271 8316 3648 8344
rect 2271 8313 2283 8316
rect 2225 8307 2283 8313
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 4212 8316 5733 8344
rect 4212 8304 4218 8316
rect 5721 8313 5733 8316
rect 5767 8313 5779 8347
rect 5721 8307 5779 8313
rect 7852 8344 7880 8375
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8386 8344 8392 8356
rect 7852 8316 8392 8344
rect 4614 8276 4620 8288
rect 4575 8248 4620 8276
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 4798 8236 4804 8288
rect 4856 8276 4862 8288
rect 7852 8276 7880 8316
rect 8386 8304 8392 8316
rect 8444 8344 8450 8356
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 8444 8316 8769 8344
rect 8444 8304 8450 8316
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 4856 8248 7880 8276
rect 4856 8236 4862 8248
rect 1104 8186 13800 8208
rect 1104 8134 3066 8186
rect 3118 8134 3130 8186
rect 3182 8134 3194 8186
rect 3246 8134 3258 8186
rect 3310 8134 3322 8186
rect 3374 8134 7298 8186
rect 7350 8134 7362 8186
rect 7414 8134 7426 8186
rect 7478 8134 7490 8186
rect 7542 8134 7554 8186
rect 7606 8134 11530 8186
rect 11582 8134 11594 8186
rect 11646 8134 11658 8186
rect 11710 8134 11722 8186
rect 11774 8134 11786 8186
rect 11838 8134 13800 8186
rect 1104 8112 13800 8134
rect 5537 8075 5595 8081
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 5718 8072 5724 8084
rect 5583 8044 5724 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 5718 8032 5724 8044
rect 5776 8072 5782 8084
rect 8205 8075 8263 8081
rect 5776 8044 7144 8072
rect 5776 8032 5782 8044
rect 7116 8004 7144 8044
rect 8205 8041 8217 8075
rect 8251 8072 8263 8075
rect 8938 8072 8944 8084
rect 8251 8044 8944 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 12066 8004 12072 8016
rect 7116 7976 12072 8004
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 2866 7936 2872 7948
rect 2827 7908 2872 7936
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 7852 7908 9321 7936
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 4157 7871 4215 7877
rect 3099 7840 3832 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 2038 7760 2044 7812
rect 2096 7800 2102 7812
rect 3602 7800 3608 7812
rect 2096 7772 3608 7800
rect 2096 7760 2102 7772
rect 3602 7760 3608 7772
rect 3660 7760 3666 7812
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3237 7735 3295 7741
rect 3237 7732 3249 7735
rect 3108 7704 3249 7732
rect 3108 7692 3114 7704
rect 3237 7701 3249 7704
rect 3283 7701 3295 7735
rect 3804 7732 3832 7840
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4706 7868 4712 7880
rect 4203 7840 4712 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4706 7828 4712 7840
rect 4764 7868 4770 7880
rect 5166 7868 5172 7880
rect 4764 7840 5172 7868
rect 4764 7828 4770 7840
rect 5166 7828 5172 7840
rect 5224 7868 5230 7880
rect 5994 7868 6000 7880
rect 5224 7840 6000 7868
rect 5224 7828 5230 7840
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 7852 7877 7880 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 11974 7868 11980 7880
rect 7837 7831 7895 7837
rect 7944 7840 11980 7868
rect 3878 7760 3884 7812
rect 3936 7800 3942 7812
rect 4402 7803 4460 7809
rect 4402 7800 4414 7803
rect 3936 7772 4414 7800
rect 3936 7760 3942 7772
rect 4402 7769 4414 7772
rect 4448 7769 4460 7803
rect 4402 7763 4460 7769
rect 5810 7760 5816 7812
rect 5868 7800 5874 7812
rect 6242 7803 6300 7809
rect 6242 7800 6254 7803
rect 5868 7772 6254 7800
rect 5868 7760 5874 7772
rect 6242 7769 6254 7772
rect 6288 7769 6300 7803
rect 6242 7763 6300 7769
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 7852 7800 7880 7831
rect 6420 7772 7880 7800
rect 6420 7760 6426 7772
rect 4614 7732 4620 7744
rect 3804 7704 4620 7732
rect 3237 7695 3295 7701
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 5592 7704 7389 7732
rect 5592 7692 5598 7704
rect 7377 7701 7389 7704
rect 7423 7732 7435 7735
rect 7944 7732 7972 7840
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 9490 7800 9496 7812
rect 9403 7772 9496 7800
rect 9490 7760 9496 7772
rect 9548 7800 9554 7812
rect 12802 7800 12808 7812
rect 9548 7772 12808 7800
rect 9548 7760 9554 7772
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 8202 7732 8208 7744
rect 7423 7704 7972 7732
rect 8163 7704 8208 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8389 7735 8447 7741
rect 8389 7701 8401 7735
rect 8435 7732 8447 7735
rect 9122 7732 9128 7744
rect 8435 7704 9128 7732
rect 8435 7701 8447 7704
rect 8389 7695 8447 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 1104 7642 13800 7664
rect 1104 7590 5182 7642
rect 5234 7590 5246 7642
rect 5298 7590 5310 7642
rect 5362 7590 5374 7642
rect 5426 7590 5438 7642
rect 5490 7590 9414 7642
rect 9466 7590 9478 7642
rect 9530 7590 9542 7642
rect 9594 7590 9606 7642
rect 9658 7590 9670 7642
rect 9722 7590 13800 7642
rect 1104 7568 13800 7590
rect 3878 7528 3884 7540
rect 3839 7500 3884 7528
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 4522 7528 4528 7540
rect 4483 7500 4528 7528
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5810 7528 5816 7540
rect 5771 7500 5816 7528
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8389 7531 8447 7537
rect 8389 7528 8401 7531
rect 8260 7500 8401 7528
rect 8260 7488 8266 7500
rect 8389 7497 8401 7500
rect 8435 7497 8447 7531
rect 8389 7491 8447 7497
rect 3602 7460 3608 7472
rect 3563 7432 3608 7460
rect 3602 7420 3608 7432
rect 3660 7420 3666 7472
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 6270 7460 6276 7472
rect 4387 7432 6276 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 6270 7420 6276 7432
rect 6328 7420 6334 7472
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 9306 7460 9312 7472
rect 8076 7432 9312 7460
rect 8076 7420 8082 7432
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2314 7352 2320 7404
rect 2372 7392 2378 7404
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2372 7364 2881 7392
rect 2372 7352 2378 7364
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 3050 7392 3056 7404
rect 3011 7364 3056 7392
rect 2869 7355 2927 7361
rect 3050 7352 3056 7364
rect 3108 7392 3114 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3108 7364 3801 7392
rect 3108 7352 3114 7364
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 4154 7392 4160 7404
rect 3927 7364 4160 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4614 7392 4620 7404
rect 4575 7364 4620 7392
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 4939 7364 5365 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 5353 7361 5365 7364
rect 5399 7392 5411 7395
rect 5534 7392 5540 7404
rect 5399 7364 5540 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 2958 7324 2964 7336
rect 2179 7296 2964 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 1964 7256 1992 7287
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 3145 7327 3203 7333
rect 3145 7293 3157 7327
rect 3191 7324 3203 7327
rect 3326 7324 3332 7336
rect 3191 7296 3332 7324
rect 3191 7293 3203 7296
rect 3145 7287 3203 7293
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 4062 7324 4068 7336
rect 3476 7296 4068 7324
rect 3476 7284 3482 7296
rect 4062 7284 4068 7296
rect 4120 7324 4126 7336
rect 4724 7324 4752 7355
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 4120 7296 4752 7324
rect 5644 7324 5672 7355
rect 6178 7352 6184 7404
rect 6236 7392 6242 7404
rect 6362 7392 6368 7404
rect 6236 7364 6368 7392
rect 6236 7352 6242 7364
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 6914 7392 6920 7404
rect 6595 7364 6920 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6914 7352 6920 7364
rect 6972 7392 6978 7404
rect 6972 7364 7696 7392
rect 6972 7352 6978 7364
rect 7668 7333 7696 7364
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8680 7401 8708 7432
rect 9306 7420 9312 7432
rect 9364 7460 9370 7472
rect 9585 7463 9643 7469
rect 9585 7460 9597 7463
rect 9364 7432 9597 7460
rect 9364 7420 9370 7432
rect 9585 7429 9597 7432
rect 9631 7429 9643 7463
rect 9585 7423 9643 7429
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7800 7364 7941 7392
rect 7800 7352 7806 7364
rect 7929 7361 7941 7364
rect 7975 7392 7987 7395
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 7975 7364 8585 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 9214 7392 9220 7404
rect 8803 7364 9220 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 9214 7352 9220 7364
rect 9272 7392 9278 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9272 7364 9413 7392
rect 9272 7352 9278 7364
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 12802 7392 12808 7404
rect 12763 7364 12808 7392
rect 9677 7355 9735 7361
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 5644 7296 6469 7324
rect 4120 7284 4126 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7293 7711 7327
rect 8846 7324 8852 7336
rect 8807 7296 8852 7324
rect 7653 7287 7711 7293
rect 7668 7256 7696 7287
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 7834 7256 7840 7268
rect 1964 7228 4200 7256
rect 7668 7228 7840 7256
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 4172 7188 4200 7228
rect 7834 7216 7840 7228
rect 7892 7256 7898 7268
rect 9692 7256 9720 7355
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 13078 7324 13084 7336
rect 13039 7296 13084 7324
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 7892 7228 9720 7256
rect 7892 7216 7898 7228
rect 4246 7188 4252 7200
rect 4159 7160 4252 7188
rect 4246 7148 4252 7160
rect 4304 7188 4310 7200
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 4304 7160 5457 7188
rect 4304 7148 4310 7160
rect 5445 7157 5457 7160
rect 5491 7157 5503 7191
rect 5445 7151 5503 7157
rect 8110 7148 8116 7200
rect 8168 7188 8174 7200
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 8168 7160 9413 7188
rect 8168 7148 8174 7160
rect 9401 7157 9413 7160
rect 9447 7157 9459 7191
rect 9401 7151 9459 7157
rect 1104 7098 13800 7120
rect 1104 7046 3066 7098
rect 3118 7046 3130 7098
rect 3182 7046 3194 7098
rect 3246 7046 3258 7098
rect 3310 7046 3322 7098
rect 3374 7046 7298 7098
rect 7350 7046 7362 7098
rect 7414 7046 7426 7098
rect 7478 7046 7490 7098
rect 7542 7046 7554 7098
rect 7606 7046 11530 7098
rect 11582 7046 11594 7098
rect 11646 7046 11658 7098
rect 11710 7046 11722 7098
rect 11774 7046 11786 7098
rect 11838 7046 13800 7098
rect 1104 7024 13800 7046
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4985 6987 5043 6993
rect 4985 6984 4997 6987
rect 4120 6956 4997 6984
rect 4120 6944 4126 6956
rect 4985 6953 4997 6956
rect 5031 6953 5043 6987
rect 4985 6947 5043 6953
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 7147 6956 8953 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4212 6888 4292 6916
rect 4212 6876 4218 6888
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3016 6820 3801 6848
rect 3016 6808 3022 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 4264 6857 4292 6888
rect 6472 6888 8064 6916
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3936 6820 4077 6848
rect 3936 6808 3942 6820
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 6472 6848 6500 6888
rect 8036 6860 8064 6888
rect 4249 6811 4307 6817
rect 6380 6820 6500 6848
rect 6380 6792 6408 6820
rect 6914 6808 6920 6860
rect 6972 6808 6978 6860
rect 8018 6848 8024 6860
rect 7979 6820 8024 6848
rect 8018 6808 8024 6820
rect 8076 6808 8082 6860
rect 8128 6857 8156 6956
rect 8941 6953 8953 6956
rect 8987 6984 8999 6987
rect 9214 6984 9220 6996
rect 8987 6956 9220 6984
rect 8987 6953 8999 6956
rect 8941 6947 8999 6953
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 1486 6780 1492 6792
rect 1447 6752 1492 6780
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 1762 6789 1768 6792
rect 1756 6743 1768 6789
rect 1820 6780 1826 6792
rect 3973 6783 4031 6789
rect 1820 6752 1856 6780
rect 1762 6740 1768 6743
rect 1820 6740 1826 6752
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 6362 6780 6368 6792
rect 4203 6752 5120 6780
rect 6275 6752 6368 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 3988 6712 4016 6743
rect 3988 6684 4568 6712
rect 4540 6656 4568 6684
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 4953 6715 5011 6721
rect 4953 6712 4965 6715
rect 4672 6684 4965 6712
rect 4672 6672 4678 6684
rect 4953 6681 4965 6684
rect 4999 6681 5011 6715
rect 4953 6675 5011 6681
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 4154 6644 4160 6656
rect 2915 6616 4160 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4580 6616 4813 6644
rect 4580 6604 4586 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 5092 6644 5120 6752
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6932 6780 6960 6808
rect 6503 6752 6960 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7892 6752 7941 6780
rect 7892 6740 7898 6752
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6780 8263 6783
rect 8386 6780 8392 6792
rect 8251 6752 8392 6780
rect 8251 6749 8263 6752
rect 8205 6743 8263 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 9030 6780 9036 6792
rect 8720 6752 9036 6780
rect 8720 6740 8726 6752
rect 9030 6740 9036 6752
rect 9088 6780 9094 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9088 6752 10333 6780
rect 9088 6740 9094 6752
rect 10321 6749 10333 6752
rect 10367 6780 10379 6783
rect 12802 6780 12808 6792
rect 10367 6752 12808 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 5166 6672 5172 6724
rect 5224 6712 5230 6724
rect 6178 6712 6184 6724
rect 5224 6684 5269 6712
rect 6139 6684 6184 6712
rect 5224 6672 5230 6684
rect 6178 6672 6184 6684
rect 6236 6672 6242 6724
rect 6917 6715 6975 6721
rect 6917 6681 6929 6715
rect 6963 6712 6975 6715
rect 7006 6712 7012 6724
rect 6963 6684 7012 6712
rect 6963 6681 6975 6684
rect 6917 6675 6975 6681
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7133 6715 7191 6721
rect 7133 6681 7145 6715
rect 7179 6712 7191 6715
rect 7179 6684 8248 6712
rect 7179 6681 7191 6684
rect 7133 6675 7191 6681
rect 5718 6644 5724 6656
rect 5092 6616 5724 6644
rect 4801 6607 4859 6613
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 6270 6644 6276 6656
rect 6328 6653 6334 6656
rect 6237 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6607 6337 6653
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7650 6644 7656 6656
rect 7331 6616 7656 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 6328 6604 6334 6607
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 7745 6647 7803 6653
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 7926 6644 7932 6656
rect 7791 6616 7932 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8220 6644 8248 6684
rect 8294 6672 8300 6724
rect 8352 6712 8358 6724
rect 10054 6715 10112 6721
rect 10054 6712 10066 6715
rect 8352 6684 10066 6712
rect 8352 6672 8358 6684
rect 10054 6681 10066 6684
rect 10100 6681 10112 6715
rect 10054 6675 10112 6681
rect 8386 6644 8392 6656
rect 8220 6616 8392 6644
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 1104 6554 13800 6576
rect 1104 6502 5182 6554
rect 5234 6502 5246 6554
rect 5298 6502 5310 6554
rect 5362 6502 5374 6554
rect 5426 6502 5438 6554
rect 5490 6502 9414 6554
rect 9466 6502 9478 6554
rect 9530 6502 9542 6554
rect 9594 6502 9606 6554
rect 9658 6502 9670 6554
rect 9722 6502 13800 6554
rect 1104 6480 13800 6502
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 5074 6440 5080 6452
rect 3476 6412 5080 6440
rect 3476 6400 3482 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 1756 6375 1814 6381
rect 1756 6341 1768 6375
rect 1802 6372 1814 6375
rect 2682 6372 2688 6384
rect 1802 6344 2688 6372
rect 1802 6341 1814 6344
rect 1756 6335 1814 6341
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 3878 6332 3884 6384
rect 3936 6372 3942 6384
rect 3936 6344 5120 6372
rect 3936 6332 3942 6344
rect 1486 6304 1492 6316
rect 1399 6276 1492 6304
rect 1486 6264 1492 6276
rect 1544 6304 1550 6316
rect 4522 6304 4528 6316
rect 1544 6276 4200 6304
rect 4483 6276 4528 6304
rect 1544 6264 1550 6276
rect 2774 6128 2780 6180
rect 2832 6168 2838 6180
rect 2869 6171 2927 6177
rect 2869 6168 2881 6171
rect 2832 6140 2881 6168
rect 2832 6128 2838 6140
rect 2869 6137 2881 6140
rect 2915 6137 2927 6171
rect 4172 6168 4200 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4982 6304 4988 6316
rect 4943 6276 4988 6304
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 5092 6313 5120 6344
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5166 6304 5172 6316
rect 5123 6276 5172 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5718 6304 5724 6316
rect 5307 6276 5724 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6328 6276 6653 6304
rect 6328 6264 6334 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 8409 6307 8467 6313
rect 8409 6273 8421 6307
rect 8455 6304 8467 6307
rect 8938 6304 8944 6316
rect 8455 6276 8944 6304
rect 8455 6273 8467 6276
rect 8409 6267 8467 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 9364 6276 9413 6304
rect 9364 6264 9370 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6236 4307 6239
rect 5000 6236 5028 6264
rect 6362 6236 6368 6248
rect 4295 6208 5028 6236
rect 6323 6208 6368 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 6362 6196 6368 6208
rect 6420 6196 6426 6248
rect 8662 6236 8668 6248
rect 8623 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9214 6236 9220 6248
rect 9171 6208 9220 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 4706 6168 4712 6180
rect 4172 6140 4712 6168
rect 2869 6131 2927 6137
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 6178 6168 6184 6180
rect 5000 6140 6184 6168
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 5000 6100 5028 6140
rect 6178 6128 6184 6140
rect 6236 6128 6242 6180
rect 6914 6168 6920 6180
rect 6472 6140 6920 6168
rect 2188 6072 5028 6100
rect 2188 6060 2194 6072
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 6472 6109 6500 6140
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 5261 6103 5319 6109
rect 5261 6100 5273 6103
rect 5132 6072 5273 6100
rect 5132 6060 5138 6072
rect 5261 6069 5273 6072
rect 5307 6069 5319 6103
rect 5261 6063 5319 6069
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 6825 6103 6883 6109
rect 6825 6069 6837 6103
rect 6871 6100 6883 6103
rect 7006 6100 7012 6112
rect 6871 6072 7012 6100
rect 6871 6069 6883 6072
rect 6825 6063 6883 6069
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7285 6103 7343 6109
rect 7285 6100 7297 6103
rect 7248 6072 7297 6100
rect 7248 6060 7254 6072
rect 7285 6069 7297 6072
rect 7331 6100 7343 6103
rect 8846 6100 8852 6112
rect 7331 6072 8852 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 1104 6010 13800 6032
rect 1104 5958 3066 6010
rect 3118 5958 3130 6010
rect 3182 5958 3194 6010
rect 3246 5958 3258 6010
rect 3310 5958 3322 6010
rect 3374 5958 7298 6010
rect 7350 5958 7362 6010
rect 7414 5958 7426 6010
rect 7478 5958 7490 6010
rect 7542 5958 7554 6010
rect 7606 5958 11530 6010
rect 11582 5958 11594 6010
rect 11646 5958 11658 6010
rect 11710 5958 11722 6010
rect 11774 5958 11786 6010
rect 11838 5958 13800 6010
rect 1104 5936 13800 5958
rect 1486 5896 1492 5908
rect 1447 5868 1492 5896
rect 1486 5856 1492 5868
rect 1544 5856 1550 5908
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 4798 5896 4804 5908
rect 3936 5868 4804 5896
rect 3936 5856 3942 5868
rect 4798 5856 4804 5868
rect 4856 5896 4862 5908
rect 4856 5868 5304 5896
rect 4856 5856 4862 5868
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 2746 5800 3801 5828
rect 2746 5760 2774 5800
rect 3789 5797 3801 5800
rect 3835 5828 3847 5831
rect 4154 5828 4160 5840
rect 3835 5800 4160 5828
rect 3835 5797 3847 5800
rect 3789 5791 3847 5797
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 5166 5828 5172 5840
rect 5092 5800 5172 5828
rect 4982 5760 4988 5772
rect 2240 5732 2774 5760
rect 2976 5732 4988 5760
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 2130 5692 2136 5704
rect 2091 5664 2136 5692
rect 1673 5655 1731 5661
rect 1688 5624 1716 5655
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 2240 5624 2268 5732
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2363 5664 2789 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2777 5661 2789 5664
rect 2823 5692 2835 5695
rect 2976 5692 3004 5732
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5092 5769 5120 5800
rect 5166 5788 5172 5800
rect 5224 5788 5230 5840
rect 5276 5769 5304 5868
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 8662 5896 8668 5908
rect 6052 5868 8668 5896
rect 6052 5856 6058 5868
rect 6932 5769 6960 5868
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 8938 5896 8944 5908
rect 8899 5868 8944 5896
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5729 5135 5763
rect 5077 5723 5135 5729
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 6917 5763 6975 5769
rect 6917 5729 6929 5763
rect 6963 5729 6975 5763
rect 6917 5723 6975 5729
rect 2823 5664 3004 5692
rect 3053 5695 3111 5701
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 3878 5692 3884 5704
rect 3099 5664 3884 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 4019 5664 5181 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 5169 5661 5181 5664
rect 5215 5661 5227 5695
rect 5169 5655 5227 5661
rect 1688 5596 2268 5624
rect 2958 5584 2964 5636
rect 3016 5624 3022 5636
rect 3418 5624 3424 5636
rect 3016 5596 3424 5624
rect 3016 5584 3022 5596
rect 3418 5584 3424 5596
rect 3476 5624 3482 5636
rect 4157 5627 4215 5633
rect 4157 5624 4169 5627
rect 3476 5596 4169 5624
rect 3476 5584 3482 5596
rect 4157 5593 4169 5596
rect 4203 5593 4215 5627
rect 4157 5587 4215 5593
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 4430 5624 4436 5636
rect 4387 5596 4436 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 5184 5624 5212 5655
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7173 5695 7231 5701
rect 7173 5692 7185 5695
rect 7064 5664 7185 5692
rect 7064 5652 7070 5664
rect 7173 5661 7185 5664
rect 7219 5661 7231 5695
rect 9122 5692 9128 5704
rect 9083 5664 9128 5692
rect 7173 5655 7231 5661
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 5718 5624 5724 5636
rect 5184 5596 5724 5624
rect 5718 5584 5724 5596
rect 5776 5584 5782 5636
rect 2866 5556 2872 5568
rect 2827 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3878 5556 3884 5568
rect 3283 5528 3884 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4801 5559 4859 5565
rect 4120 5528 4165 5556
rect 4120 5516 4126 5528
rect 4801 5525 4813 5559
rect 4847 5556 4859 5559
rect 4890 5556 4896 5568
rect 4847 5528 4896 5556
rect 4847 5525 4859 5528
rect 4801 5519 4859 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8386 5556 8392 5568
rect 8343 5528 8392 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8386 5516 8392 5528
rect 8444 5556 8450 5568
rect 9214 5556 9220 5568
rect 8444 5528 9220 5556
rect 8444 5516 8450 5528
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 1104 5466 13800 5488
rect 1104 5414 5182 5466
rect 5234 5414 5246 5466
rect 5298 5414 5310 5466
rect 5362 5414 5374 5466
rect 5426 5414 5438 5466
rect 5490 5414 9414 5466
rect 9466 5414 9478 5466
rect 9530 5414 9542 5466
rect 9594 5414 9606 5466
rect 9658 5414 9670 5466
rect 9722 5414 13800 5466
rect 1104 5392 13800 5414
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 8294 5352 8300 5364
rect 8067 5324 8300 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 4706 5284 4712 5296
rect 4356 5256 4712 5284
rect 4356 5228 4384 5256
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 3053 5219 3111 5225
rect 3053 5216 3065 5219
rect 3016 5188 3065 5216
rect 3016 5176 3022 5188
rect 3053 5185 3065 5188
rect 3099 5216 3111 5219
rect 4062 5216 4068 5228
rect 3099 5188 4068 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4338 5216 4344 5228
rect 4251 5188 4344 5216
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4614 5225 4620 5228
rect 4608 5179 4620 5225
rect 4672 5216 4678 5228
rect 7926 5216 7932 5228
rect 4672 5188 4708 5216
rect 7887 5188 7932 5216
rect 4614 5176 4620 5179
rect 4672 5176 4678 5188
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 8110 5216 8116 5228
rect 8071 5188 8116 5216
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3329 5151 3387 5157
rect 3329 5148 3341 5151
rect 2924 5120 3341 5148
rect 2924 5108 2930 5120
rect 3329 5117 3341 5120
rect 3375 5148 3387 5151
rect 3786 5148 3792 5160
rect 3375 5120 3792 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 5718 5080 5724 5092
rect 5631 5052 5724 5080
rect 5718 5040 5724 5052
rect 5776 5080 5782 5092
rect 12618 5080 12624 5092
rect 5776 5052 12624 5080
rect 5776 5040 5782 5052
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 1104 4922 13800 4944
rect 1104 4870 3066 4922
rect 3118 4870 3130 4922
rect 3182 4870 3194 4922
rect 3246 4870 3258 4922
rect 3310 4870 3322 4922
rect 3374 4870 7298 4922
rect 7350 4870 7362 4922
rect 7414 4870 7426 4922
rect 7478 4870 7490 4922
rect 7542 4870 7554 4922
rect 7606 4870 11530 4922
rect 11582 4870 11594 4922
rect 11646 4870 11658 4922
rect 11710 4870 11722 4922
rect 11774 4870 11786 4922
rect 11838 4870 13800 4922
rect 1104 4848 13800 4870
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4672 4780 4905 4808
rect 4672 4768 4678 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 4893 4771 4951 4777
rect 4982 4672 4988 4684
rect 4264 4644 4988 4672
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4264 4613 4292 4644
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3936 4576 3985 4604
rect 3936 4564 3942 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4890 4604 4896 4616
rect 4851 4576 4896 4604
rect 4433 4567 4491 4573
rect 3804 4536 3832 4564
rect 4448 4536 4476 4567
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 3804 4508 4476 4536
rect 3786 4468 3792 4480
rect 3747 4440 3792 4468
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 1104 4378 13800 4400
rect 1104 4326 5182 4378
rect 5234 4326 5246 4378
rect 5298 4326 5310 4378
rect 5362 4326 5374 4378
rect 5426 4326 5438 4378
rect 5490 4326 9414 4378
rect 9466 4326 9478 4378
rect 9530 4326 9542 4378
rect 9594 4326 9606 4378
rect 9658 4326 9670 4378
rect 9722 4326 13800 4378
rect 1104 4304 13800 4326
rect 3636 4199 3694 4205
rect 3636 4165 3648 4199
rect 3682 4196 3694 4199
rect 3786 4196 3792 4208
rect 3682 4168 3792 4196
rect 3682 4165 3694 4168
rect 3636 4159 3694 4165
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 4338 4128 4344 4140
rect 3927 4100 4344 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 2501 3927 2559 3933
rect 2501 3893 2513 3927
rect 2547 3924 2559 3927
rect 2958 3924 2964 3936
rect 2547 3896 2964 3924
rect 2547 3893 2559 3896
rect 2501 3887 2559 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 1104 3834 13800 3856
rect 1104 3782 3066 3834
rect 3118 3782 3130 3834
rect 3182 3782 3194 3834
rect 3246 3782 3258 3834
rect 3310 3782 3322 3834
rect 3374 3782 7298 3834
rect 7350 3782 7362 3834
rect 7414 3782 7426 3834
rect 7478 3782 7490 3834
rect 7542 3782 7554 3834
rect 7606 3782 11530 3834
rect 11582 3782 11594 3834
rect 11646 3782 11658 3834
rect 11710 3782 11722 3834
rect 11774 3782 11786 3834
rect 11838 3782 13800 3834
rect 1104 3760 13800 3782
rect 12802 3584 12808 3596
rect 12763 3556 12808 3584
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 13078 3516 13084 3528
rect 13039 3488 13084 3516
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 1104 3290 13800 3312
rect 1104 3238 5182 3290
rect 5234 3238 5246 3290
rect 5298 3238 5310 3290
rect 5362 3238 5374 3290
rect 5426 3238 5438 3290
rect 5490 3238 9414 3290
rect 9466 3238 9478 3290
rect 9530 3238 9542 3290
rect 9594 3238 9606 3290
rect 9658 3238 9670 3290
rect 9722 3238 13800 3290
rect 1104 3216 13800 3238
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2958 3040 2964 3052
rect 1719 3012 2964 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 1486 2836 1492 2848
rect 1447 2808 1492 2836
rect 1486 2796 1492 2808
rect 1544 2796 1550 2848
rect 1104 2746 13800 2768
rect 1104 2694 3066 2746
rect 3118 2694 3130 2746
rect 3182 2694 3194 2746
rect 3246 2694 3258 2746
rect 3310 2694 3322 2746
rect 3374 2694 7298 2746
rect 7350 2694 7362 2746
rect 7414 2694 7426 2746
rect 7478 2694 7490 2746
rect 7542 2694 7554 2746
rect 7606 2694 11530 2746
rect 11582 2694 11594 2746
rect 11646 2694 11658 2746
rect 11710 2694 11722 2746
rect 11774 2694 11786 2746
rect 11838 2694 13800 2746
rect 1104 2672 13800 2694
rect 11974 2524 11980 2576
rect 12032 2564 12038 2576
rect 12989 2567 13047 2573
rect 12989 2564 13001 2567
rect 12032 2536 13001 2564
rect 12032 2524 12038 2536
rect 12989 2533 13001 2536
rect 13035 2533 13047 2567
rect 12989 2527 13047 2533
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2958 2428 2964 2440
rect 2919 2400 2964 2428
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7190 2428 7196 2440
rect 6687 2400 7196 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9214 2428 9220 2440
rect 9171 2400 9220 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 12066 2428 12072 2440
rect 12027 2400 12072 2428
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12492 2400 12817 2428
rect 12492 2388 12498 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1489 2295 1547 2301
rect 1489 2292 1501 2295
rect 72 2264 1501 2292
rect 72 2252 78 2264
rect 1489 2261 1501 2264
rect 1535 2261 1547 2295
rect 1489 2255 1547 2261
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 2777 2295 2835 2301
rect 2777 2292 2789 2295
rect 2648 2264 2789 2292
rect 2648 2252 2654 2264
rect 2777 2261 2789 2264
rect 2823 2261 2835 2295
rect 2777 2255 2835 2261
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 5868 2264 6469 2292
rect 5868 2252 5874 2264
rect 6457 2261 6469 2264
rect 6503 2261 6515 2295
rect 6457 2255 6515 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 12250 2292 12256 2304
rect 12211 2264 12256 2292
rect 9309 2255 9367 2261
rect 12250 2252 12256 2264
rect 12308 2252 12314 2304
rect 1104 2202 13800 2224
rect 1104 2150 5182 2202
rect 5234 2150 5246 2202
rect 5298 2150 5310 2202
rect 5362 2150 5374 2202
rect 5426 2150 5438 2202
rect 5490 2150 9414 2202
rect 9466 2150 9478 2202
rect 9530 2150 9542 2202
rect 9594 2150 9606 2202
rect 9658 2150 9670 2202
rect 9722 2150 13800 2202
rect 1104 2128 13800 2150
<< via1 >>
rect 3066 14662 3118 14714
rect 3130 14662 3182 14714
rect 3194 14662 3246 14714
rect 3258 14662 3310 14714
rect 3322 14662 3374 14714
rect 7298 14662 7350 14714
rect 7362 14662 7414 14714
rect 7426 14662 7478 14714
rect 7490 14662 7542 14714
rect 7554 14662 7606 14714
rect 11530 14662 11582 14714
rect 11594 14662 11646 14714
rect 11658 14662 11710 14714
rect 11722 14662 11774 14714
rect 11786 14662 11838 14714
rect 1492 14603 1544 14612
rect 1492 14569 1501 14603
rect 1501 14569 1535 14603
rect 1535 14569 1544 14603
rect 1492 14560 1544 14569
rect 2780 14603 2832 14612
rect 2780 14569 2789 14603
rect 2789 14569 2823 14603
rect 2823 14569 2832 14603
rect 2780 14560 2832 14569
rect 5816 14560 5868 14612
rect 9036 14560 9088 14612
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 14832 14560 14884 14612
rect 4160 14356 4212 14408
rect 5908 14356 5960 14408
rect 9312 14356 9364 14408
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 12440 14356 12492 14408
rect 4804 14288 4856 14340
rect 5182 14118 5234 14170
rect 5246 14118 5298 14170
rect 5310 14118 5362 14170
rect 5374 14118 5426 14170
rect 5438 14118 5490 14170
rect 9414 14118 9466 14170
rect 9478 14118 9530 14170
rect 9542 14118 9594 14170
rect 9606 14118 9658 14170
rect 9670 14118 9722 14170
rect 10324 13880 10376 13932
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 3066 13574 3118 13626
rect 3130 13574 3182 13626
rect 3194 13574 3246 13626
rect 3258 13574 3310 13626
rect 3322 13574 3374 13626
rect 7298 13574 7350 13626
rect 7362 13574 7414 13626
rect 7426 13574 7478 13626
rect 7490 13574 7542 13626
rect 7554 13574 7606 13626
rect 11530 13574 11582 13626
rect 11594 13574 11646 13626
rect 11658 13574 11710 13626
rect 11722 13574 11774 13626
rect 11786 13574 11838 13626
rect 7196 13268 7248 13320
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 5182 13030 5234 13082
rect 5246 13030 5298 13082
rect 5310 13030 5362 13082
rect 5374 13030 5426 13082
rect 5438 13030 5490 13082
rect 9414 13030 9466 13082
rect 9478 13030 9530 13082
rect 9542 13030 9594 13082
rect 9606 13030 9658 13082
rect 9670 13030 9722 13082
rect 3066 12486 3118 12538
rect 3130 12486 3182 12538
rect 3194 12486 3246 12538
rect 3258 12486 3310 12538
rect 3322 12486 3374 12538
rect 7298 12486 7350 12538
rect 7362 12486 7414 12538
rect 7426 12486 7478 12538
rect 7490 12486 7542 12538
rect 7554 12486 7606 12538
rect 11530 12486 11582 12538
rect 11594 12486 11646 12538
rect 11658 12486 11710 12538
rect 11722 12486 11774 12538
rect 11786 12486 11838 12538
rect 5182 11942 5234 11994
rect 5246 11942 5298 11994
rect 5310 11942 5362 11994
rect 5374 11942 5426 11994
rect 5438 11942 5490 11994
rect 9414 11942 9466 11994
rect 9478 11942 9530 11994
rect 9542 11942 9594 11994
rect 9606 11942 9658 11994
rect 9670 11942 9722 11994
rect 6368 11636 6420 11688
rect 6920 11611 6972 11620
rect 6920 11577 6929 11611
rect 6929 11577 6963 11611
rect 6963 11577 6972 11611
rect 6920 11568 6972 11577
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 3066 11398 3118 11450
rect 3130 11398 3182 11450
rect 3194 11398 3246 11450
rect 3258 11398 3310 11450
rect 3322 11398 3374 11450
rect 7298 11398 7350 11450
rect 7362 11398 7414 11450
rect 7426 11398 7478 11450
rect 7490 11398 7542 11450
rect 7554 11398 7606 11450
rect 11530 11398 11582 11450
rect 11594 11398 11646 11450
rect 11658 11398 11710 11450
rect 11722 11398 11774 11450
rect 11786 11398 11838 11450
rect 7196 11296 7248 11348
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 5632 11160 5684 11212
rect 8116 11203 8168 11212
rect 8116 11169 8125 11203
rect 8125 11169 8159 11203
rect 8159 11169 8168 11203
rect 8116 11160 8168 11169
rect 9864 11160 9916 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 7932 11135 7984 11144
rect 5080 11024 5132 11076
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 6460 11024 6512 11076
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 2412 10956 2464 11008
rect 4620 10999 4672 11008
rect 4620 10965 4629 10999
rect 4629 10965 4663 10999
rect 4663 10965 4672 10999
rect 4620 10956 4672 10965
rect 8208 10956 8260 11008
rect 5182 10854 5234 10906
rect 5246 10854 5298 10906
rect 5310 10854 5362 10906
rect 5374 10854 5426 10906
rect 5438 10854 5490 10906
rect 9414 10854 9466 10906
rect 9478 10854 9530 10906
rect 9542 10854 9594 10906
rect 9606 10854 9658 10906
rect 9670 10854 9722 10906
rect 4160 10752 4212 10804
rect 5632 10795 5684 10804
rect 5632 10761 5641 10795
rect 5641 10761 5675 10795
rect 5675 10761 5684 10795
rect 5632 10752 5684 10761
rect 7104 10752 7156 10804
rect 7196 10752 7248 10804
rect 2872 10684 2924 10736
rect 2044 10659 2096 10668
rect 2044 10625 2078 10659
rect 2078 10625 2096 10659
rect 6552 10684 6604 10736
rect 2044 10616 2096 10625
rect 3792 10616 3844 10668
rect 5080 10616 5132 10668
rect 7380 10616 7432 10668
rect 5908 10548 5960 10600
rect 10324 10616 10376 10668
rect 12624 10616 12676 10668
rect 8208 10548 8260 10600
rect 8760 10548 8812 10600
rect 3424 10412 3476 10464
rect 12440 10548 12492 10600
rect 9864 10523 9916 10532
rect 9864 10489 9873 10523
rect 9873 10489 9907 10523
rect 9907 10489 9916 10523
rect 9864 10480 9916 10489
rect 7932 10412 7984 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 3066 10310 3118 10362
rect 3130 10310 3182 10362
rect 3194 10310 3246 10362
rect 3258 10310 3310 10362
rect 3322 10310 3374 10362
rect 7298 10310 7350 10362
rect 7362 10310 7414 10362
rect 7426 10310 7478 10362
rect 7490 10310 7542 10362
rect 7554 10310 7606 10362
rect 11530 10310 11582 10362
rect 11594 10310 11646 10362
rect 11658 10310 11710 10362
rect 11722 10310 11774 10362
rect 11786 10310 11838 10362
rect 2044 10208 2096 10260
rect 2596 10208 2648 10260
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 5172 10208 5224 10260
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 6460 10251 6512 10260
rect 6460 10217 6469 10251
rect 6469 10217 6503 10251
rect 6503 10217 6512 10251
rect 6460 10208 6512 10217
rect 6920 10208 6972 10260
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 7196 10072 7248 10124
rect 7932 10072 7984 10124
rect 2412 10004 2464 10013
rect 3424 10004 3476 10056
rect 4620 10004 4672 10056
rect 7012 10004 7064 10056
rect 7656 10004 7708 10056
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 9036 10004 9088 10056
rect 2688 9936 2740 9988
rect 4896 9936 4948 9988
rect 7840 9936 7892 9988
rect 9220 9979 9272 9988
rect 9220 9945 9254 9979
rect 9254 9945 9272 9979
rect 9220 9936 9272 9945
rect 7748 9868 7800 9920
rect 9036 9868 9088 9920
rect 5182 9766 5234 9818
rect 5246 9766 5298 9818
rect 5310 9766 5362 9818
rect 5374 9766 5426 9818
rect 5438 9766 5490 9818
rect 9414 9766 9466 9818
rect 9478 9766 9530 9818
rect 9542 9766 9594 9818
rect 9606 9766 9658 9818
rect 9670 9766 9722 9818
rect 3792 9707 3844 9716
rect 3792 9673 3801 9707
rect 3801 9673 3835 9707
rect 3835 9673 3844 9707
rect 3792 9664 3844 9673
rect 4160 9664 4212 9716
rect 2136 9528 2188 9580
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 1676 9324 1728 9376
rect 3792 9324 3844 9376
rect 4988 9460 5040 9512
rect 6552 9596 6604 9648
rect 5908 9528 5960 9580
rect 6920 9596 6972 9648
rect 8024 9596 8076 9648
rect 8116 9596 8168 9648
rect 8392 9528 8444 9580
rect 9588 9571 9640 9580
rect 9588 9537 9622 9571
rect 9622 9537 9640 9571
rect 6368 9503 6420 9512
rect 6368 9469 6377 9503
rect 6377 9469 6411 9503
rect 6411 9469 6420 9503
rect 6368 9460 6420 9469
rect 6552 9503 6604 9512
rect 6552 9469 6561 9503
rect 6561 9469 6595 9503
rect 6595 9469 6604 9503
rect 6552 9460 6604 9469
rect 7104 9460 7156 9512
rect 7564 9460 7616 9512
rect 8116 9460 8168 9512
rect 8208 9460 8260 9512
rect 9588 9528 9640 9537
rect 9128 9460 9180 9512
rect 7932 9392 7984 9444
rect 6368 9324 6420 9376
rect 8024 9324 8076 9376
rect 8208 9324 8260 9376
rect 8944 9324 8996 9376
rect 12440 9324 12492 9376
rect 3066 9222 3118 9274
rect 3130 9222 3182 9274
rect 3194 9222 3246 9274
rect 3258 9222 3310 9274
rect 3322 9222 3374 9274
rect 7298 9222 7350 9274
rect 7362 9222 7414 9274
rect 7426 9222 7478 9274
rect 7490 9222 7542 9274
rect 7554 9222 7606 9274
rect 11530 9222 11582 9274
rect 11594 9222 11646 9274
rect 11658 9222 11710 9274
rect 11722 9222 11774 9274
rect 11786 9222 11838 9274
rect 1676 9120 1728 9172
rect 4620 9120 4672 9172
rect 4896 9120 4948 9172
rect 8760 9120 8812 9172
rect 9220 9163 9272 9172
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 9588 9120 9640 9172
rect 6920 8984 6972 9036
rect 7932 9027 7984 9036
rect 7932 8993 7941 9027
rect 7941 8993 7975 9027
rect 7975 8993 7984 9027
rect 7932 8984 7984 8993
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 7656 8916 7708 8968
rect 8392 8916 8444 8968
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 9036 8959 9088 8968
rect 9036 8925 9045 8959
rect 9045 8925 9079 8959
rect 9079 8925 9088 8959
rect 9036 8916 9088 8925
rect 10048 8916 10100 8968
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 2412 8891 2464 8900
rect 2412 8857 2421 8891
rect 2421 8857 2455 8891
rect 2455 8857 2464 8891
rect 2412 8848 2464 8857
rect 2596 8891 2648 8900
rect 2596 8857 2621 8891
rect 2621 8857 2648 8891
rect 3792 8891 3844 8900
rect 2596 8848 2648 8857
rect 3792 8857 3801 8891
rect 3801 8857 3835 8891
rect 3835 8857 3844 8891
rect 3792 8848 3844 8857
rect 4528 8848 4580 8900
rect 4804 8891 4856 8900
rect 4804 8857 4813 8891
rect 4813 8857 4847 8891
rect 4847 8857 4856 8891
rect 4804 8848 4856 8857
rect 1768 8823 1820 8832
rect 1768 8789 1783 8823
rect 1783 8789 1817 8823
rect 1817 8789 1820 8823
rect 1768 8780 1820 8789
rect 2872 8780 2924 8832
rect 3332 8780 3384 8832
rect 4252 8780 4304 8832
rect 7748 8848 7800 8900
rect 8300 8848 8352 8900
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 5182 8678 5234 8730
rect 5246 8678 5298 8730
rect 5310 8678 5362 8730
rect 5374 8678 5426 8730
rect 5438 8678 5490 8730
rect 9414 8678 9466 8730
rect 9478 8678 9530 8730
rect 9542 8678 9594 8730
rect 9606 8678 9658 8730
rect 9670 8678 9722 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 2044 8508 2096 8560
rect 2688 8508 2740 8560
rect 1768 8440 1820 8492
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 4160 8440 4212 8492
rect 7840 8508 7892 8560
rect 3792 8372 3844 8424
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 7748 8440 7800 8492
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 8392 8440 8444 8492
rect 9496 8440 9548 8492
rect 6276 8372 6328 8424
rect 8024 8415 8076 8424
rect 4160 8304 4212 8356
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 4804 8236 4856 8288
rect 8392 8304 8444 8356
rect 3066 8134 3118 8186
rect 3130 8134 3182 8186
rect 3194 8134 3246 8186
rect 3258 8134 3310 8186
rect 3322 8134 3374 8186
rect 7298 8134 7350 8186
rect 7362 8134 7414 8186
rect 7426 8134 7478 8186
rect 7490 8134 7542 8186
rect 7554 8134 7606 8186
rect 11530 8134 11582 8186
rect 11594 8134 11646 8186
rect 11658 8134 11710 8186
rect 11722 8134 11774 8186
rect 11786 8134 11838 8186
rect 5724 8032 5776 8084
rect 8944 8032 8996 8084
rect 12072 7964 12124 8016
rect 2872 7939 2924 7948
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 2872 7896 2924 7905
rect 2044 7760 2096 7812
rect 3608 7760 3660 7812
rect 3056 7692 3108 7744
rect 4712 7828 4764 7880
rect 5172 7828 5224 7880
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6000 7828 6052 7837
rect 3884 7760 3936 7812
rect 5816 7760 5868 7812
rect 6368 7760 6420 7812
rect 4620 7692 4672 7744
rect 5540 7692 5592 7744
rect 11980 7828 12032 7880
rect 9496 7803 9548 7812
rect 9496 7769 9505 7803
rect 9505 7769 9539 7803
rect 9539 7769 9548 7803
rect 9496 7760 9548 7769
rect 12808 7760 12860 7812
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 9128 7692 9180 7744
rect 5182 7590 5234 7642
rect 5246 7590 5298 7642
rect 5310 7590 5362 7642
rect 5374 7590 5426 7642
rect 5438 7590 5490 7642
rect 9414 7590 9466 7642
rect 9478 7590 9530 7642
rect 9542 7590 9594 7642
rect 9606 7590 9658 7642
rect 9670 7590 9722 7642
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 8208 7488 8260 7540
rect 3608 7463 3660 7472
rect 3608 7429 3617 7463
rect 3617 7429 3651 7463
rect 3651 7429 3660 7463
rect 3608 7420 3660 7429
rect 6276 7420 6328 7472
rect 8024 7420 8076 7472
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2320 7352 2372 7404
rect 3056 7395 3108 7404
rect 3056 7361 3065 7395
rect 3065 7361 3099 7395
rect 3099 7361 3108 7395
rect 3056 7352 3108 7361
rect 4160 7352 4212 7404
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 2964 7284 3016 7336
rect 3332 7284 3384 7336
rect 3424 7284 3476 7336
rect 4068 7284 4120 7336
rect 5540 7352 5592 7404
rect 6184 7352 6236 7404
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 6920 7352 6972 7404
rect 7748 7352 7800 7404
rect 9312 7420 9364 7472
rect 9220 7352 9272 7404
rect 12808 7395 12860 7404
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 7840 7216 7892 7268
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 13084 7327 13136 7336
rect 13084 7293 13093 7327
rect 13093 7293 13127 7327
rect 13127 7293 13136 7327
rect 13084 7284 13136 7293
rect 4252 7148 4304 7200
rect 8116 7148 8168 7200
rect 3066 7046 3118 7098
rect 3130 7046 3182 7098
rect 3194 7046 3246 7098
rect 3258 7046 3310 7098
rect 3322 7046 3374 7098
rect 7298 7046 7350 7098
rect 7362 7046 7414 7098
rect 7426 7046 7478 7098
rect 7490 7046 7542 7098
rect 7554 7046 7606 7098
rect 11530 7046 11582 7098
rect 11594 7046 11646 7098
rect 11658 7046 11710 7098
rect 11722 7046 11774 7098
rect 11786 7046 11838 7098
rect 4068 6944 4120 6996
rect 4160 6876 4212 6928
rect 2964 6808 3016 6860
rect 3884 6808 3936 6860
rect 6920 6808 6972 6860
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 8024 6808 8076 6817
rect 9220 6944 9272 6996
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 1768 6783 1820 6792
rect 1768 6749 1802 6783
rect 1802 6749 1820 6783
rect 1768 6740 1820 6749
rect 6368 6783 6420 6792
rect 4620 6672 4672 6724
rect 4160 6604 4212 6656
rect 4528 6604 4580 6656
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 7840 6740 7892 6792
rect 8392 6740 8444 6792
rect 8668 6740 8720 6792
rect 9036 6740 9088 6792
rect 12808 6740 12860 6792
rect 5172 6715 5224 6724
rect 5172 6681 5181 6715
rect 5181 6681 5215 6715
rect 5215 6681 5224 6715
rect 6184 6715 6236 6724
rect 5172 6672 5224 6681
rect 6184 6681 6193 6715
rect 6193 6681 6227 6715
rect 6227 6681 6236 6715
rect 6184 6672 6236 6681
rect 7012 6672 7064 6724
rect 5724 6604 5776 6656
rect 6276 6647 6328 6656
rect 6276 6613 6291 6647
rect 6291 6613 6325 6647
rect 6325 6613 6328 6647
rect 6276 6604 6328 6613
rect 7656 6604 7708 6656
rect 7932 6604 7984 6656
rect 8300 6672 8352 6724
rect 8392 6604 8444 6656
rect 5182 6502 5234 6554
rect 5246 6502 5298 6554
rect 5310 6502 5362 6554
rect 5374 6502 5426 6554
rect 5438 6502 5490 6554
rect 9414 6502 9466 6554
rect 9478 6502 9530 6554
rect 9542 6502 9594 6554
rect 9606 6502 9658 6554
rect 9670 6502 9722 6554
rect 3424 6400 3476 6452
rect 5080 6400 5132 6452
rect 2688 6332 2740 6384
rect 3884 6332 3936 6384
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 4528 6307 4580 6316
rect 1492 6264 1544 6273
rect 2780 6128 2832 6180
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5172 6264 5224 6316
rect 5724 6264 5776 6316
rect 6276 6264 6328 6316
rect 8944 6264 8996 6316
rect 9312 6264 9364 6316
rect 6368 6239 6420 6248
rect 6368 6205 6377 6239
rect 6377 6205 6411 6239
rect 6411 6205 6420 6239
rect 6368 6196 6420 6205
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 9220 6196 9272 6248
rect 4712 6128 4764 6180
rect 2136 6060 2188 6112
rect 6184 6128 6236 6180
rect 5080 6060 5132 6112
rect 6920 6128 6972 6180
rect 7012 6060 7064 6112
rect 7196 6060 7248 6112
rect 8852 6060 8904 6112
rect 3066 5958 3118 6010
rect 3130 5958 3182 6010
rect 3194 5958 3246 6010
rect 3258 5958 3310 6010
rect 3322 5958 3374 6010
rect 7298 5958 7350 6010
rect 7362 5958 7414 6010
rect 7426 5958 7478 6010
rect 7490 5958 7542 6010
rect 7554 5958 7606 6010
rect 11530 5958 11582 6010
rect 11594 5958 11646 6010
rect 11658 5958 11710 6010
rect 11722 5958 11774 6010
rect 11786 5958 11838 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 3884 5856 3936 5908
rect 4804 5856 4856 5908
rect 4160 5788 4212 5840
rect 4988 5763 5040 5772
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 4988 5729 4997 5763
rect 4997 5729 5031 5763
rect 5031 5729 5040 5763
rect 4988 5720 5040 5729
rect 5172 5788 5224 5840
rect 6000 5856 6052 5908
rect 8668 5856 8720 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 3884 5652 3936 5704
rect 2964 5584 3016 5636
rect 3424 5584 3476 5636
rect 4436 5584 4488 5636
rect 7012 5652 7064 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 5724 5584 5776 5636
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 3884 5516 3936 5568
rect 4068 5559 4120 5568
rect 4068 5525 4077 5559
rect 4077 5525 4111 5559
rect 4111 5525 4120 5559
rect 4068 5516 4120 5525
rect 4896 5516 4948 5568
rect 8392 5516 8444 5568
rect 9220 5516 9272 5568
rect 5182 5414 5234 5466
rect 5246 5414 5298 5466
rect 5310 5414 5362 5466
rect 5374 5414 5426 5466
rect 5438 5414 5490 5466
rect 9414 5414 9466 5466
rect 9478 5414 9530 5466
rect 9542 5414 9594 5466
rect 9606 5414 9658 5466
rect 9670 5414 9722 5466
rect 8300 5312 8352 5364
rect 4712 5244 4764 5296
rect 2964 5176 3016 5228
rect 4068 5176 4120 5228
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 4620 5219 4672 5228
rect 4620 5185 4654 5219
rect 4654 5185 4672 5219
rect 7932 5219 7984 5228
rect 4620 5176 4672 5185
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 2872 5108 2924 5160
rect 3792 5108 3844 5160
rect 5724 5083 5776 5092
rect 5724 5049 5733 5083
rect 5733 5049 5767 5083
rect 5767 5049 5776 5083
rect 5724 5040 5776 5049
rect 12624 5040 12676 5092
rect 3066 4870 3118 4922
rect 3130 4870 3182 4922
rect 3194 4870 3246 4922
rect 3258 4870 3310 4922
rect 3322 4870 3374 4922
rect 7298 4870 7350 4922
rect 7362 4870 7414 4922
rect 7426 4870 7478 4922
rect 7490 4870 7542 4922
rect 7554 4870 7606 4922
rect 11530 4870 11582 4922
rect 11594 4870 11646 4922
rect 11658 4870 11710 4922
rect 11722 4870 11774 4922
rect 11786 4870 11838 4922
rect 4620 4768 4672 4820
rect 3792 4564 3844 4616
rect 3884 4564 3936 4616
rect 4988 4632 5040 4684
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 5182 4326 5234 4378
rect 5246 4326 5298 4378
rect 5310 4326 5362 4378
rect 5374 4326 5426 4378
rect 5438 4326 5490 4378
rect 9414 4326 9466 4378
rect 9478 4326 9530 4378
rect 9542 4326 9594 4378
rect 9606 4326 9658 4378
rect 9670 4326 9722 4378
rect 3792 4156 3844 4208
rect 4344 4088 4396 4140
rect 2964 3884 3016 3936
rect 3066 3782 3118 3834
rect 3130 3782 3182 3834
rect 3194 3782 3246 3834
rect 3258 3782 3310 3834
rect 3322 3782 3374 3834
rect 7298 3782 7350 3834
rect 7362 3782 7414 3834
rect 7426 3782 7478 3834
rect 7490 3782 7542 3834
rect 7554 3782 7606 3834
rect 11530 3782 11582 3834
rect 11594 3782 11646 3834
rect 11658 3782 11710 3834
rect 11722 3782 11774 3834
rect 11786 3782 11838 3834
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 5182 3238 5234 3290
rect 5246 3238 5298 3290
rect 5310 3238 5362 3290
rect 5374 3238 5426 3290
rect 5438 3238 5490 3290
rect 9414 3238 9466 3290
rect 9478 3238 9530 3290
rect 9542 3238 9594 3290
rect 9606 3238 9658 3290
rect 9670 3238 9722 3290
rect 2964 3000 3016 3052
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 3066 2694 3118 2746
rect 3130 2694 3182 2746
rect 3194 2694 3246 2746
rect 3258 2694 3310 2746
rect 3322 2694 3374 2746
rect 7298 2694 7350 2746
rect 7362 2694 7414 2746
rect 7426 2694 7478 2746
rect 7490 2694 7542 2746
rect 7554 2694 7606 2746
rect 11530 2694 11582 2746
rect 11594 2694 11646 2746
rect 11658 2694 11710 2746
rect 11722 2694 11774 2746
rect 11786 2694 11838 2746
rect 11980 2524 12032 2576
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 7196 2388 7248 2440
rect 9220 2388 9272 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12440 2388 12492 2440
rect 20 2252 72 2304
rect 2596 2252 2648 2304
rect 5816 2252 5868 2304
rect 9036 2252 9088 2304
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 5182 2150 5234 2202
rect 5246 2150 5298 2202
rect 5310 2150 5362 2202
rect 5374 2150 5426 2202
rect 5438 2150 5490 2202
rect 9414 2150 9466 2202
rect 9478 2150 9530 2202
rect 9542 2150 9594 2202
rect 9606 2150 9658 2202
rect 9670 2150 9722 2202
<< metal2 >>
rect 1490 16416 1546 16425
rect 1490 16351 1546 16360
rect 1504 14618 1532 16351
rect 2594 16325 2650 17125
rect 5814 16325 5870 17125
rect 9034 16325 9090 17125
rect 12254 16325 12310 17125
rect 14830 16325 14886 17125
rect 2608 15178 2636 16325
rect 2608 15150 2820 15178
rect 2792 14618 2820 15150
rect 3066 14716 3374 14736
rect 3066 14714 3072 14716
rect 3128 14714 3152 14716
rect 3208 14714 3232 14716
rect 3288 14714 3312 14716
rect 3368 14714 3374 14716
rect 3128 14662 3130 14714
rect 3310 14662 3312 14714
rect 3066 14660 3072 14662
rect 3128 14660 3152 14662
rect 3208 14660 3232 14662
rect 3288 14660 3312 14662
rect 3368 14660 3374 14662
rect 3066 14640 3374 14660
rect 5828 14618 5856 16325
rect 7298 14716 7606 14736
rect 7298 14714 7304 14716
rect 7360 14714 7384 14716
rect 7440 14714 7464 14716
rect 7520 14714 7544 14716
rect 7600 14714 7606 14716
rect 7360 14662 7362 14714
rect 7542 14662 7544 14714
rect 7298 14660 7304 14662
rect 7360 14660 7384 14662
rect 7440 14660 7464 14662
rect 7520 14660 7544 14662
rect 7600 14660 7606 14662
rect 7298 14640 7606 14660
rect 9048 14618 9076 16325
rect 11530 14716 11838 14736
rect 11530 14714 11536 14716
rect 11592 14714 11616 14716
rect 11672 14714 11696 14716
rect 11752 14714 11776 14716
rect 11832 14714 11838 14716
rect 11592 14662 11594 14714
rect 11774 14662 11776 14714
rect 11530 14660 11536 14662
rect 11592 14660 11616 14662
rect 11672 14660 11696 14662
rect 11752 14660 11776 14662
rect 11832 14660 11838 14662
rect 11530 14640 11838 14660
rect 12268 14618 12296 16325
rect 14844 14618 14872 16325
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 3066 13628 3374 13648
rect 3066 13626 3072 13628
rect 3128 13626 3152 13628
rect 3208 13626 3232 13628
rect 3288 13626 3312 13628
rect 3368 13626 3374 13628
rect 3128 13574 3130 13626
rect 3310 13574 3312 13626
rect 3066 13572 3072 13574
rect 3128 13572 3152 13574
rect 3208 13572 3232 13574
rect 3288 13572 3312 13574
rect 3368 13572 3374 13574
rect 3066 13552 3374 13572
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 13025 1532 13126
rect 1490 13016 1546 13025
rect 1490 12951 1546 12960
rect 3066 12540 3374 12560
rect 3066 12538 3072 12540
rect 3128 12538 3152 12540
rect 3208 12538 3232 12540
rect 3288 12538 3312 12540
rect 3368 12538 3374 12540
rect 3128 12486 3130 12538
rect 3310 12486 3312 12538
rect 3066 12484 3072 12486
rect 3128 12484 3152 12486
rect 3208 12484 3232 12486
rect 3288 12484 3312 12486
rect 3368 12484 3374 12486
rect 3066 12464 3374 12484
rect 3066 11452 3374 11472
rect 3066 11450 3072 11452
rect 3128 11450 3152 11452
rect 3208 11450 3232 11452
rect 3288 11450 3312 11452
rect 3368 11450 3374 11452
rect 3128 11398 3130 11450
rect 3310 11398 3312 11450
rect 3066 11396 3072 11398
rect 3128 11396 3152 11398
rect 3208 11396 3232 11398
rect 3288 11396 3312 11398
rect 3368 11396 3374 11398
rect 3066 11376 3374 11396
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 9625 1440 11086
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 10266 2084 10610
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2424 10062 2452 10950
rect 4172 10810 4200 14350
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4816 11218 4844 14282
rect 5182 14172 5490 14192
rect 5182 14170 5188 14172
rect 5244 14170 5268 14172
rect 5324 14170 5348 14172
rect 5404 14170 5428 14172
rect 5484 14170 5490 14172
rect 5244 14118 5246 14170
rect 5426 14118 5428 14170
rect 5182 14116 5188 14118
rect 5244 14116 5268 14118
rect 5324 14116 5348 14118
rect 5404 14116 5428 14118
rect 5484 14116 5490 14118
rect 5182 14096 5490 14116
rect 5182 13084 5490 13104
rect 5182 13082 5188 13084
rect 5244 13082 5268 13084
rect 5324 13082 5348 13084
rect 5404 13082 5428 13084
rect 5484 13082 5490 13084
rect 5244 13030 5246 13082
rect 5426 13030 5428 13082
rect 5182 13028 5188 13030
rect 5244 13028 5268 13030
rect 5324 13028 5348 13030
rect 5404 13028 5428 13030
rect 5484 13028 5490 13030
rect 5182 13008 5490 13028
rect 5182 11996 5490 12016
rect 5182 11994 5188 11996
rect 5244 11994 5268 11996
rect 5324 11994 5348 11996
rect 5404 11994 5428 11996
rect 5484 11994 5490 11996
rect 5244 11942 5246 11994
rect 5426 11942 5428 11994
rect 5182 11940 5188 11942
rect 5244 11940 5268 11942
rect 5324 11940 5348 11942
rect 5404 11940 5428 11942
rect 5484 11940 5490 11942
rect 5182 11920 5490 11940
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 9178 1716 9318
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1688 8906 1716 9114
rect 1676 8900 1728 8906
rect 1676 8842 1728 8848
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1504 6322 1532 6734
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1490 6216 1546 6225
rect 1490 6151 1546 6160
rect 1504 5914 1532 6151
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1492 2848 1544 2854
rect 1490 2816 1492 2825
rect 1544 2816 1546 2825
rect 1490 2751 1546 2760
rect 1688 2446 1716 8842
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8498 1808 8774
rect 2148 8634 2176 9522
rect 2424 8906 2452 9998
rect 2608 8906 2636 10202
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2700 8566 2728 9930
rect 2884 9586 2912 10678
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3066 10364 3374 10384
rect 3066 10362 3072 10364
rect 3128 10362 3152 10364
rect 3208 10362 3232 10364
rect 3288 10362 3312 10364
rect 3368 10362 3374 10364
rect 3128 10310 3130 10362
rect 3310 10310 3312 10362
rect 3066 10308 3072 10310
rect 3128 10308 3152 10310
rect 3208 10308 3232 10310
rect 3288 10308 3312 10310
rect 3368 10308 3374 10310
rect 3066 10288 3374 10308
rect 3436 10062 3464 10406
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3804 9722 3832 10610
rect 4172 9722 4200 10746
rect 4632 10062 4660 10950
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4908 9994 4936 11086
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3066 9276 3374 9296
rect 3066 9274 3072 9276
rect 3128 9274 3152 9276
rect 3208 9274 3232 9276
rect 3288 9274 3312 9276
rect 3368 9274 3374 9276
rect 3128 9222 3130 9274
rect 3310 9222 3312 9274
rect 3066 9220 3072 9222
rect 3128 9220 3152 9222
rect 3208 9220 3232 9222
rect 3288 9220 3312 9222
rect 3368 9220 3374 9222
rect 3066 9200 3374 9220
rect 3804 8906 3832 9318
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 2044 8560 2096 8566
rect 2044 8502 2096 8508
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 2056 7818 2084 8502
rect 2884 7954 2912 8774
rect 3344 8498 3372 8774
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 8378 3372 8434
rect 3804 8430 3832 8842
rect 4172 8498 4200 9658
rect 4908 9178 4936 9930
rect 5000 9518 5028 11086
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 10674 5120 11018
rect 5182 10908 5490 10928
rect 5182 10906 5188 10908
rect 5244 10906 5268 10908
rect 5324 10906 5348 10908
rect 5404 10906 5428 10908
rect 5484 10906 5490 10908
rect 5244 10854 5246 10906
rect 5426 10854 5428 10906
rect 5182 10852 5188 10854
rect 5244 10852 5268 10854
rect 5324 10852 5348 10854
rect 5404 10852 5428 10854
rect 5484 10852 5490 10854
rect 5182 10832 5490 10852
rect 5644 10810 5672 11154
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10248 5120 10610
rect 5920 10606 5948 14350
rect 7298 13628 7606 13648
rect 7298 13626 7304 13628
rect 7360 13626 7384 13628
rect 7440 13626 7464 13628
rect 7520 13626 7544 13628
rect 7600 13626 7606 13628
rect 7360 13574 7362 13626
rect 7542 13574 7544 13626
rect 7298 13572 7304 13574
rect 7360 13572 7384 13574
rect 7440 13572 7464 13574
rect 7520 13572 7544 13574
rect 7600 13572 7606 13574
rect 7298 13552 7606 13572
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5920 10266 5948 10542
rect 5172 10260 5224 10266
rect 5092 10220 5172 10248
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3792 8424 3844 8430
rect 3344 8350 3464 8378
rect 3792 8366 3844 8372
rect 3066 8188 3374 8208
rect 3066 8186 3072 8188
rect 3128 8186 3152 8188
rect 3208 8186 3232 8188
rect 3288 8186 3312 8188
rect 3368 8186 3374 8188
rect 3128 8134 3130 8186
rect 3310 8134 3312 8186
rect 3066 8132 3072 8134
rect 3128 8132 3152 8134
rect 3208 8132 3232 8134
rect 3288 8132 3312 8134
rect 3368 8132 3374 8134
rect 3066 8112 3374 8132
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2044 7812 2096 7818
rect 2044 7754 2096 7760
rect 2056 7410 2084 7754
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3068 7410 3096 7686
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1780 6798 1808 7142
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5710 2176 6054
rect 2332 5914 2360 7346
rect 3436 7342 3464 8350
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3620 7478 3648 7754
rect 3896 7546 3924 7754
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 4172 7410 4200 8298
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2700 6390 2728 7142
rect 2976 6866 3004 7278
rect 3344 7188 3372 7278
rect 3344 7160 3464 7188
rect 3066 7100 3374 7120
rect 3066 7098 3072 7100
rect 3128 7098 3152 7100
rect 3208 7098 3232 7100
rect 3288 7098 3312 7100
rect 3368 7098 3374 7100
rect 3128 7046 3130 7098
rect 3310 7046 3312 7098
rect 3066 7044 3072 7046
rect 3128 7044 3152 7046
rect 3208 7044 3232 7046
rect 3288 7044 3312 7046
rect 3368 7044 3374 7046
rect 3066 7024 3374 7044
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 3436 6458 3464 7160
rect 4080 7002 4108 7278
rect 4264 7206 4292 8774
rect 4540 7546 4568 8842
rect 4632 8294 4660 9114
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4816 8294 4844 8842
rect 5092 8548 5120 10220
rect 5172 10202 5224 10208
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5182 9820 5490 9840
rect 5182 9818 5188 9820
rect 5244 9818 5268 9820
rect 5324 9818 5348 9820
rect 5404 9818 5428 9820
rect 5484 9818 5490 9820
rect 5244 9766 5246 9818
rect 5426 9766 5428 9818
rect 5182 9764 5188 9766
rect 5244 9764 5268 9766
rect 5324 9764 5348 9766
rect 5404 9764 5428 9766
rect 5484 9764 5490 9766
rect 5182 9744 5490 9764
rect 5920 9586 5948 10202
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 6380 9518 6408 11630
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6472 10266 6500 11018
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6564 9654 6592 10678
rect 6932 10266 6960 11562
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7024 10062 7052 11494
rect 7208 11354 7236 13262
rect 7298 12540 7606 12560
rect 7298 12538 7304 12540
rect 7360 12538 7384 12540
rect 7440 12538 7464 12540
rect 7520 12538 7544 12540
rect 7600 12538 7606 12540
rect 7360 12486 7362 12538
rect 7542 12486 7544 12538
rect 7298 12484 7304 12486
rect 7360 12484 7384 12486
rect 7440 12484 7464 12486
rect 7520 12484 7544 12486
rect 7600 12484 7606 12486
rect 7298 12464 7606 12484
rect 7298 11452 7606 11472
rect 7298 11450 7304 11452
rect 7360 11450 7384 11452
rect 7440 11450 7464 11452
rect 7520 11450 7544 11452
rect 7600 11450 7606 11452
rect 7360 11398 7362 11450
rect 7542 11398 7544 11450
rect 7298 11396 7304 11398
rect 7360 11396 7384 11398
rect 7440 11396 7464 11398
rect 7520 11396 7544 11398
rect 7600 11396 7606 11398
rect 7298 11376 7606 11396
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7208 10810 7236 11290
rect 8036 11218 8156 11234
rect 8036 11212 8168 11218
rect 8036 11206 8116 11212
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6564 9518 6592 9590
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 5182 8732 5490 8752
rect 5182 8730 5188 8732
rect 5244 8730 5268 8732
rect 5324 8730 5348 8732
rect 5404 8730 5428 8732
rect 5484 8730 5490 8732
rect 5244 8678 5246 8730
rect 5426 8678 5428 8730
rect 5182 8676 5188 8678
rect 5244 8676 5268 8678
rect 5324 8676 5348 8678
rect 5404 8676 5428 8678
rect 5484 8676 5490 8678
rect 5182 8656 5490 8676
rect 5092 8520 5212 8548
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4632 7750 4660 8230
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2792 5658 2820 6122
rect 3066 6012 3374 6032
rect 3066 6010 3072 6012
rect 3128 6010 3152 6012
rect 3208 6010 3232 6012
rect 3288 6010 3312 6012
rect 3368 6010 3374 6012
rect 3128 5958 3130 6010
rect 3310 5958 3312 6010
rect 3066 5956 3072 5958
rect 3128 5956 3152 5958
rect 3208 5956 3232 5958
rect 3288 5956 3312 5958
rect 3368 5956 3374 5958
rect 3066 5936 3374 5956
rect 2792 5642 3004 5658
rect 3436 5642 3464 6394
rect 3896 6390 3924 6802
rect 4172 6662 4200 6870
rect 4540 6746 4568 7482
rect 4632 7410 4660 7686
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4448 6718 4568 6746
rect 4632 6730 4660 7346
rect 4620 6724 4672 6730
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 3884 6384 3936 6390
rect 3804 6344 3884 6372
rect 2792 5636 3016 5642
rect 2792 5630 2964 5636
rect 2792 2774 2820 5630
rect 2964 5578 3016 5584
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5166 2912 5510
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2976 3942 3004 5170
rect 3804 5166 3832 6344
rect 3884 6326 3936 6332
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3896 5710 3924 5850
rect 4172 5846 4200 6598
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 4448 5642 4476 6718
rect 4620 6666 4672 6672
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6322 4568 6598
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4724 6186 4752 7822
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3066 4924 3374 4944
rect 3066 4922 3072 4924
rect 3128 4922 3152 4924
rect 3208 4922 3232 4924
rect 3288 4922 3312 4924
rect 3368 4922 3374 4924
rect 3128 4870 3130 4922
rect 3310 4870 3312 4922
rect 3066 4868 3072 4870
rect 3128 4868 3152 4870
rect 3208 4868 3232 4870
rect 3288 4868 3312 4870
rect 3368 4868 3374 4870
rect 3066 4848 3374 4868
rect 3804 4622 3832 5102
rect 3896 4622 3924 5510
rect 4080 5234 4108 5510
rect 4724 5302 4752 6122
rect 4816 5914 4844 8230
rect 5184 7886 5212 8520
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5736 8090 5764 8434
rect 6288 8430 6316 8910
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5182 7644 5490 7664
rect 5182 7642 5188 7644
rect 5244 7642 5268 7644
rect 5324 7642 5348 7644
rect 5404 7642 5428 7644
rect 5484 7642 5490 7644
rect 5244 7590 5246 7642
rect 5426 7590 5428 7642
rect 5182 7588 5188 7590
rect 5244 7588 5268 7590
rect 5324 7588 5348 7590
rect 5404 7588 5428 7590
rect 5484 7588 5490 7590
rect 5182 7568 5490 7588
rect 5552 7410 5580 7686
rect 5828 7546 5856 7754
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5092 6730 5212 6746
rect 5092 6724 5224 6730
rect 5092 6718 5172 6724
rect 5092 6458 5120 6718
rect 5172 6666 5224 6672
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5182 6556 5490 6576
rect 5182 6554 5188 6556
rect 5244 6554 5268 6556
rect 5324 6554 5348 6556
rect 5404 6554 5428 6556
rect 5484 6554 5490 6556
rect 5244 6502 5246 6554
rect 5426 6502 5428 6554
rect 5182 6500 5188 6502
rect 5244 6500 5268 6502
rect 5324 6500 5348 6502
rect 5404 6500 5428 6502
rect 5484 6500 5490 6502
rect 5182 6480 5490 6500
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5736 6322 5764 6598
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5000 5778 5028 6258
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 4214 3832 4422
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 4356 4146 4384 5170
rect 4632 4826 4660 5170
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4908 4622 4936 5510
rect 5000 4690 5028 5714
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5092 4622 5120 6054
rect 5184 5846 5212 6258
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 5736 5642 5764 6258
rect 6012 5914 6040 7822
rect 6288 7478 6316 8366
rect 6380 7818 6408 9318
rect 6932 9042 6960 9590
rect 7116 9518 7144 10746
rect 7208 10130 7236 10746
rect 7380 10668 7432 10674
rect 7432 10628 7788 10656
rect 7380 10610 7432 10616
rect 7298 10364 7606 10384
rect 7298 10362 7304 10364
rect 7360 10362 7384 10364
rect 7440 10362 7464 10364
rect 7520 10362 7544 10364
rect 7600 10362 7606 10364
rect 7360 10310 7362 10362
rect 7542 10310 7544 10362
rect 7298 10308 7304 10310
rect 7360 10308 7384 10310
rect 7440 10308 7464 10310
rect 7520 10308 7544 10310
rect 7600 10308 7606 10310
rect 7298 10288 7606 10308
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7564 9512 7616 9518
rect 7668 9466 7696 9998
rect 7760 9926 7788 10628
rect 7944 10470 7972 11086
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10130 7972 10406
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7616 9460 7696 9466
rect 7564 9454 7696 9460
rect 7576 9438 7696 9454
rect 7298 9276 7606 9296
rect 7298 9274 7304 9276
rect 7360 9274 7384 9276
rect 7440 9274 7464 9276
rect 7520 9274 7544 9276
rect 7600 9274 7606 9276
rect 7360 9222 7362 9274
rect 7542 9222 7544 9274
rect 7298 9220 7304 9222
rect 7360 9220 7384 9222
rect 7440 9220 7464 9222
rect 7520 9220 7544 9222
rect 7600 9220 7606 9222
rect 7298 9200 7606 9220
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 7668 8974 7696 9438
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7298 8188 7606 8208
rect 7298 8186 7304 8188
rect 7360 8186 7384 8188
rect 7440 8186 7464 8188
rect 7520 8186 7544 8188
rect 7600 8186 7606 8188
rect 7360 8134 7362 8186
rect 7542 8134 7544 8186
rect 7298 8132 7304 8134
rect 7360 8132 7384 8134
rect 7440 8132 7464 8134
rect 7520 8132 7544 8134
rect 7600 8132 7606 8134
rect 7298 8112 7606 8132
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6380 7410 6408 7754
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6196 6730 6224 7346
rect 6932 6866 6960 7346
rect 7298 7100 7606 7120
rect 7298 7098 7304 7100
rect 7360 7098 7384 7100
rect 7440 7098 7464 7100
rect 7520 7098 7544 7100
rect 7600 7098 7606 7100
rect 7360 7046 7362 7098
rect 7542 7046 7544 7098
rect 7298 7044 7304 7046
rect 7360 7044 7384 7046
rect 7440 7044 7464 7046
rect 7520 7044 7544 7046
rect 7600 7044 7606 7046
rect 7298 7024 7606 7044
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6196 6186 6224 6666
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6322 6316 6598
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6380 6254 6408 6734
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6932 6186 6960 6802
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7024 6610 7052 6666
rect 7668 6662 7696 8910
rect 7760 8906 7788 9862
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7760 8498 7788 8842
rect 7852 8838 7880 9930
rect 7944 9450 7972 10066
rect 8036 9654 8064 11206
rect 8116 11154 8168 11160
rect 8208 11144 8260 11150
rect 8128 11092 8208 11098
rect 8128 11086 8260 11092
rect 8128 11070 8248 11086
rect 8128 9654 8156 11070
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10606 8248 10950
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8220 10062 8248 10542
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7944 9042 7972 9386
rect 8036 9382 8064 9590
rect 8128 9518 8156 9590
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8566 7880 8774
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 7410 7788 8434
rect 8036 8430 8064 9318
rect 8128 8498 8156 9454
rect 8220 9382 8248 9454
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8404 8974 8432 9522
rect 8772 9178 8800 10542
rect 9036 10056 9088 10062
rect 9088 10016 9168 10044
rect 9036 9998 9088 10004
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8956 8974 8984 9318
rect 9048 8974 9076 9862
rect 9140 9518 9168 10016
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8312 8634 8340 8842
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8404 8498 8432 8910
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7546 8248 7686
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7852 6798 7880 7210
rect 8036 6866 8064 7414
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7656 6656 7708 6662
rect 7024 6582 7236 6610
rect 7656 6598 7708 6604
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7208 6118 7236 6582
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 7024 5710 7052 6054
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5182 5468 5490 5488
rect 5182 5466 5188 5468
rect 5244 5466 5268 5468
rect 5324 5466 5348 5468
rect 5404 5466 5428 5468
rect 5484 5466 5490 5468
rect 5244 5414 5246 5466
rect 5426 5414 5428 5466
rect 5182 5412 5188 5414
rect 5244 5412 5268 5414
rect 5324 5412 5348 5414
rect 5404 5412 5428 5414
rect 5484 5412 5490 5414
rect 5182 5392 5490 5412
rect 5736 5098 5764 5578
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5182 4380 5490 4400
rect 5182 4378 5188 4380
rect 5244 4378 5268 4380
rect 5324 4378 5348 4380
rect 5404 4378 5428 4380
rect 5484 4378 5490 4380
rect 5244 4326 5246 4378
rect 5426 4326 5428 4378
rect 5182 4324 5188 4326
rect 5244 4324 5268 4326
rect 5324 4324 5348 4326
rect 5404 4324 5428 4326
rect 5484 4324 5490 4326
rect 5182 4304 5490 4324
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2976 3058 3004 3878
rect 3066 3836 3374 3856
rect 3066 3834 3072 3836
rect 3128 3834 3152 3836
rect 3208 3834 3232 3836
rect 3288 3834 3312 3836
rect 3368 3834 3374 3836
rect 3128 3782 3130 3834
rect 3310 3782 3312 3834
rect 3066 3780 3072 3782
rect 3128 3780 3152 3782
rect 3208 3780 3232 3782
rect 3288 3780 3312 3782
rect 3368 3780 3374 3782
rect 3066 3760 3374 3780
rect 5182 3292 5490 3312
rect 5182 3290 5188 3292
rect 5244 3290 5268 3292
rect 5324 3290 5348 3292
rect 5404 3290 5428 3292
rect 5484 3290 5490 3292
rect 5244 3238 5246 3290
rect 5426 3238 5428 3290
rect 5182 3236 5188 3238
rect 5244 3236 5268 3238
rect 5324 3236 5348 3238
rect 5404 3236 5428 3238
rect 5484 3236 5490 3238
rect 5182 3216 5490 3236
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2792 2746 3004 2774
rect 2976 2446 3004 2746
rect 3066 2748 3374 2768
rect 3066 2746 3072 2748
rect 3128 2746 3152 2748
rect 3208 2746 3232 2748
rect 3288 2746 3312 2748
rect 3368 2746 3374 2748
rect 3128 2694 3130 2746
rect 3310 2694 3312 2746
rect 3066 2692 3072 2694
rect 3128 2692 3152 2694
rect 3208 2692 3232 2694
rect 3288 2692 3312 2694
rect 3368 2692 3374 2694
rect 3066 2672 3374 2692
rect 7208 2446 7236 6054
rect 7298 6012 7606 6032
rect 7298 6010 7304 6012
rect 7360 6010 7384 6012
rect 7440 6010 7464 6012
rect 7520 6010 7544 6012
rect 7600 6010 7606 6012
rect 7360 5958 7362 6010
rect 7542 5958 7544 6010
rect 7298 5956 7304 5958
rect 7360 5956 7384 5958
rect 7440 5956 7464 5958
rect 7520 5956 7544 5958
rect 7600 5956 7606 5958
rect 7298 5936 7606 5956
rect 7944 5234 7972 6598
rect 8128 5234 8156 7142
rect 8404 6798 8432 8298
rect 8956 8090 8984 8910
rect 9140 8786 9168 9454
rect 9232 9178 9260 9930
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9048 8758 9168 8786
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8312 5370 8340 6666
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 5574 8432 6598
rect 8680 6254 8708 6734
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8680 5914 8708 6190
rect 8864 6118 8892 7278
rect 9048 6798 9076 8758
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8956 5914 8984 6258
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9140 5710 9168 7686
rect 9324 7562 9352 14350
rect 9414 14172 9722 14192
rect 9414 14170 9420 14172
rect 9476 14170 9500 14172
rect 9556 14170 9580 14172
rect 9636 14170 9660 14172
rect 9716 14170 9722 14172
rect 9476 14118 9478 14170
rect 9658 14118 9660 14170
rect 9414 14116 9420 14118
rect 9476 14116 9500 14118
rect 9556 14116 9580 14118
rect 9636 14116 9660 14118
rect 9716 14116 9722 14118
rect 9414 14096 9722 14116
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 9414 13084 9722 13104
rect 9414 13082 9420 13084
rect 9476 13082 9500 13084
rect 9556 13082 9580 13084
rect 9636 13082 9660 13084
rect 9716 13082 9722 13084
rect 9476 13030 9478 13082
rect 9658 13030 9660 13082
rect 9414 13028 9420 13030
rect 9476 13028 9500 13030
rect 9556 13028 9580 13030
rect 9636 13028 9660 13030
rect 9716 13028 9722 13030
rect 9414 13008 9722 13028
rect 9414 11996 9722 12016
rect 9414 11994 9420 11996
rect 9476 11994 9500 11996
rect 9556 11994 9580 11996
rect 9636 11994 9660 11996
rect 9716 11994 9722 11996
rect 9476 11942 9478 11994
rect 9658 11942 9660 11994
rect 9414 11940 9420 11942
rect 9476 11940 9500 11942
rect 9556 11940 9580 11942
rect 9636 11940 9660 11942
rect 9716 11940 9722 11942
rect 9414 11920 9722 11940
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9414 10908 9722 10928
rect 9414 10906 9420 10908
rect 9476 10906 9500 10908
rect 9556 10906 9580 10908
rect 9636 10906 9660 10908
rect 9716 10906 9722 10908
rect 9476 10854 9478 10906
rect 9658 10854 9660 10906
rect 9414 10852 9420 10854
rect 9476 10852 9500 10854
rect 9556 10852 9580 10854
rect 9636 10852 9660 10854
rect 9716 10852 9722 10854
rect 9414 10832 9722 10852
rect 9876 10538 9904 11154
rect 10336 10674 10364 13874
rect 11530 13628 11838 13648
rect 11530 13626 11536 13628
rect 11592 13626 11616 13628
rect 11672 13626 11696 13628
rect 11752 13626 11776 13628
rect 11832 13626 11838 13628
rect 11592 13574 11594 13626
rect 11774 13574 11776 13626
rect 11530 13572 11536 13574
rect 11592 13572 11616 13574
rect 11672 13572 11696 13574
rect 11752 13572 11776 13574
rect 11832 13572 11838 13574
rect 11530 13552 11838 13572
rect 11530 12540 11838 12560
rect 11530 12538 11536 12540
rect 11592 12538 11616 12540
rect 11672 12538 11696 12540
rect 11752 12538 11776 12540
rect 11832 12538 11838 12540
rect 11592 12486 11594 12538
rect 11774 12486 11776 12538
rect 11530 12484 11536 12486
rect 11592 12484 11616 12486
rect 11672 12484 11696 12486
rect 11752 12484 11776 12486
rect 11832 12484 11838 12486
rect 11530 12464 11838 12484
rect 12084 12434 12112 14350
rect 11992 12406 12112 12434
rect 11530 11452 11838 11472
rect 11530 11450 11536 11452
rect 11592 11450 11616 11452
rect 11672 11450 11696 11452
rect 11752 11450 11776 11452
rect 11832 11450 11838 11452
rect 11592 11398 11594 11450
rect 11774 11398 11776 11450
rect 11530 11396 11536 11398
rect 11592 11396 11616 11398
rect 11672 11396 11696 11398
rect 11752 11396 11776 11398
rect 11832 11396 11838 11398
rect 11530 11376 11838 11396
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9414 9820 9722 9840
rect 9414 9818 9420 9820
rect 9476 9818 9500 9820
rect 9556 9818 9580 9820
rect 9636 9818 9660 9820
rect 9716 9818 9722 9820
rect 9476 9766 9478 9818
rect 9658 9766 9660 9818
rect 9414 9764 9420 9766
rect 9476 9764 9500 9766
rect 9556 9764 9580 9766
rect 9636 9764 9660 9766
rect 9716 9764 9722 9766
rect 9414 9744 9722 9764
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9178 9628 9522
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 10060 8974 10088 10406
rect 10336 10266 10364 10610
rect 11530 10364 11838 10384
rect 11530 10362 11536 10364
rect 11592 10362 11616 10364
rect 11672 10362 11696 10364
rect 11752 10362 11776 10364
rect 11832 10362 11838 10364
rect 11592 10310 11594 10362
rect 11774 10310 11776 10362
rect 11530 10308 11536 10310
rect 11592 10308 11616 10310
rect 11672 10308 11696 10310
rect 11752 10308 11776 10310
rect 11832 10308 11838 10310
rect 11530 10288 11838 10308
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 11530 9276 11838 9296
rect 11530 9274 11536 9276
rect 11592 9274 11616 9276
rect 11672 9274 11696 9276
rect 11752 9274 11776 9276
rect 11832 9274 11838 9276
rect 11592 9222 11594 9274
rect 11774 9222 11776 9274
rect 11530 9220 11536 9222
rect 11592 9220 11616 9222
rect 11672 9220 11696 9222
rect 11752 9220 11776 9222
rect 11832 9220 11838 9222
rect 11530 9200 11838 9220
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9414 8732 9722 8752
rect 9414 8730 9420 8732
rect 9476 8730 9500 8732
rect 9556 8730 9580 8732
rect 9636 8730 9660 8732
rect 9716 8730 9722 8732
rect 9476 8678 9478 8730
rect 9658 8678 9660 8730
rect 9414 8676 9420 8678
rect 9476 8676 9500 8678
rect 9556 8676 9580 8678
rect 9636 8676 9660 8678
rect 9716 8676 9722 8678
rect 9414 8656 9722 8676
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9508 7818 9536 8434
rect 11530 8188 11838 8208
rect 11530 8186 11536 8188
rect 11592 8186 11616 8188
rect 11672 8186 11696 8188
rect 11752 8186 11776 8188
rect 11832 8186 11838 8188
rect 11592 8134 11594 8186
rect 11774 8134 11776 8186
rect 11530 8132 11536 8134
rect 11592 8132 11616 8134
rect 11672 8132 11696 8134
rect 11752 8132 11776 8134
rect 11832 8132 11838 8134
rect 11530 8112 11838 8132
rect 11992 7886 12020 12406
rect 12452 10606 12480 14350
rect 12992 13728 13044 13734
rect 12990 13696 12992 13705
rect 13044 13696 13046 13705
rect 12990 13631 13046 13640
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9414 7644 9722 7664
rect 9414 7642 9420 7644
rect 9476 7642 9500 7644
rect 9556 7642 9580 7644
rect 9636 7642 9660 7644
rect 9716 7642 9722 7644
rect 9476 7590 9478 7642
rect 9658 7590 9660 7642
rect 9414 7588 9420 7590
rect 9476 7588 9500 7590
rect 9556 7588 9580 7590
rect 9636 7588 9660 7590
rect 9716 7588 9722 7590
rect 9414 7568 9722 7588
rect 9232 7534 9352 7562
rect 9232 7410 9260 7534
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9232 7002 9260 7346
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9324 6322 9352 7414
rect 11530 7100 11838 7120
rect 11530 7098 11536 7100
rect 11592 7098 11616 7100
rect 11672 7098 11696 7100
rect 11752 7098 11776 7100
rect 11832 7098 11838 7100
rect 11592 7046 11594 7098
rect 11774 7046 11776 7098
rect 11530 7044 11536 7046
rect 11592 7044 11616 7046
rect 11672 7044 11696 7046
rect 11752 7044 11776 7046
rect 11832 7044 11838 7046
rect 11530 7024 11838 7044
rect 9414 6556 9722 6576
rect 9414 6554 9420 6556
rect 9476 6554 9500 6556
rect 9556 6554 9580 6556
rect 9636 6554 9660 6556
rect 9716 6554 9722 6556
rect 9476 6502 9478 6554
rect 9658 6502 9660 6554
rect 9414 6500 9420 6502
rect 9476 6500 9500 6502
rect 9556 6500 9580 6502
rect 9636 6500 9660 6502
rect 9716 6500 9722 6502
rect 9414 6480 9722 6500
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9232 5574 9260 6190
rect 11530 6012 11838 6032
rect 11530 6010 11536 6012
rect 11592 6010 11616 6012
rect 11672 6010 11696 6012
rect 11752 6010 11776 6012
rect 11832 6010 11838 6012
rect 11592 5958 11594 6010
rect 11774 5958 11776 6010
rect 11530 5956 11536 5958
rect 11592 5956 11616 5958
rect 11672 5956 11696 5958
rect 11752 5956 11776 5958
rect 11832 5956 11838 5958
rect 11530 5936 11838 5956
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7298 4924 7606 4944
rect 7298 4922 7304 4924
rect 7360 4922 7384 4924
rect 7440 4922 7464 4924
rect 7520 4922 7544 4924
rect 7600 4922 7606 4924
rect 7360 4870 7362 4922
rect 7542 4870 7544 4922
rect 7298 4868 7304 4870
rect 7360 4868 7384 4870
rect 7440 4868 7464 4870
rect 7520 4868 7544 4870
rect 7600 4868 7606 4870
rect 7298 4848 7606 4868
rect 7298 3836 7606 3856
rect 7298 3834 7304 3836
rect 7360 3834 7384 3836
rect 7440 3834 7464 3836
rect 7520 3834 7544 3836
rect 7600 3834 7606 3836
rect 7360 3782 7362 3834
rect 7542 3782 7544 3834
rect 7298 3780 7304 3782
rect 7360 3780 7384 3782
rect 7440 3780 7464 3782
rect 7520 3780 7544 3782
rect 7600 3780 7606 3782
rect 7298 3760 7606 3780
rect 7298 2748 7606 2768
rect 7298 2746 7304 2748
rect 7360 2746 7384 2748
rect 7440 2746 7464 2748
rect 7520 2746 7544 2748
rect 7600 2746 7606 2748
rect 7360 2694 7362 2746
rect 7542 2694 7544 2746
rect 7298 2692 7304 2694
rect 7360 2692 7384 2694
rect 7440 2692 7464 2694
rect 7520 2692 7544 2694
rect 7600 2692 7606 2694
rect 7298 2672 7606 2692
rect 9232 2446 9260 5510
rect 9414 5468 9722 5488
rect 9414 5466 9420 5468
rect 9476 5466 9500 5468
rect 9556 5466 9580 5468
rect 9636 5466 9660 5468
rect 9716 5466 9722 5468
rect 9476 5414 9478 5466
rect 9658 5414 9660 5466
rect 9414 5412 9420 5414
rect 9476 5412 9500 5414
rect 9556 5412 9580 5414
rect 9636 5412 9660 5414
rect 9716 5412 9722 5414
rect 9414 5392 9722 5412
rect 11530 4924 11838 4944
rect 11530 4922 11536 4924
rect 11592 4922 11616 4924
rect 11672 4922 11696 4924
rect 11752 4922 11776 4924
rect 11832 4922 11838 4924
rect 11592 4870 11594 4922
rect 11774 4870 11776 4922
rect 11530 4868 11536 4870
rect 11592 4868 11616 4870
rect 11672 4868 11696 4870
rect 11752 4868 11776 4870
rect 11832 4868 11838 4870
rect 11530 4848 11838 4868
rect 9414 4380 9722 4400
rect 9414 4378 9420 4380
rect 9476 4378 9500 4380
rect 9556 4378 9580 4380
rect 9636 4378 9660 4380
rect 9716 4378 9722 4380
rect 9476 4326 9478 4378
rect 9658 4326 9660 4378
rect 9414 4324 9420 4326
rect 9476 4324 9500 4326
rect 9556 4324 9580 4326
rect 9636 4324 9660 4326
rect 9716 4324 9722 4326
rect 9414 4304 9722 4324
rect 11530 3836 11838 3856
rect 11530 3834 11536 3836
rect 11592 3834 11616 3836
rect 11672 3834 11696 3836
rect 11752 3834 11776 3836
rect 11832 3834 11838 3836
rect 11592 3782 11594 3834
rect 11774 3782 11776 3834
rect 11530 3780 11536 3782
rect 11592 3780 11616 3782
rect 11672 3780 11696 3782
rect 11752 3780 11776 3782
rect 11832 3780 11838 3782
rect 11530 3760 11838 3780
rect 9414 3292 9722 3312
rect 9414 3290 9420 3292
rect 9476 3290 9500 3292
rect 9556 3290 9580 3292
rect 9636 3290 9660 3292
rect 9716 3290 9722 3292
rect 9476 3238 9478 3290
rect 9658 3238 9660 3290
rect 9414 3236 9420 3238
rect 9476 3236 9500 3238
rect 9556 3236 9580 3238
rect 9636 3236 9660 3238
rect 9716 3236 9722 3238
rect 9414 3216 9722 3236
rect 11530 2748 11838 2768
rect 11530 2746 11536 2748
rect 11592 2746 11616 2748
rect 11672 2746 11696 2748
rect 11752 2746 11776 2748
rect 11832 2746 11838 2748
rect 11592 2694 11594 2746
rect 11774 2694 11776 2746
rect 11530 2692 11536 2694
rect 11592 2692 11616 2694
rect 11672 2692 11696 2694
rect 11752 2692 11776 2694
rect 11832 2692 11838 2694
rect 11530 2672 11838 2692
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 32 800 60 2246
rect 2608 800 2636 2246
rect 5182 2204 5490 2224
rect 5182 2202 5188 2204
rect 5244 2202 5268 2204
rect 5324 2202 5348 2204
rect 5404 2202 5428 2204
rect 5484 2202 5490 2204
rect 5244 2150 5246 2202
rect 5426 2150 5428 2202
rect 5182 2148 5188 2150
rect 5244 2148 5268 2150
rect 5324 2148 5348 2150
rect 5404 2148 5428 2150
rect 5484 2148 5490 2150
rect 5182 2128 5490 2148
rect 5828 800 5856 2246
rect 9048 800 9076 2246
rect 9414 2204 9722 2224
rect 9414 2202 9420 2204
rect 9476 2202 9500 2204
rect 9556 2202 9580 2204
rect 9636 2202 9660 2204
rect 9716 2202 9722 2204
rect 9476 2150 9478 2202
rect 9658 2150 9660 2202
rect 9414 2148 9420 2150
rect 9476 2148 9500 2150
rect 9556 2148 9580 2150
rect 9636 2148 9660 2150
rect 9716 2148 9722 2150
rect 9414 2128 9722 2148
rect 18 0 74 800
rect 2594 0 2650 800
rect 5814 0 5870 800
rect 9034 0 9090 800
rect 11992 105 12020 2518
rect 12084 2446 12112 7958
rect 12452 2446 12480 9318
rect 12636 5098 12664 10610
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10305 13032 10406
rect 12990 10296 13046 10305
rect 12990 10231 13046 10240
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12820 7410 12848 7754
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13096 6905 13124 7278
rect 13082 6896 13138 6905
rect 13082 6831 13138 6840
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12820 3602 12848 6734
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 13084 3528 13136 3534
rect 13082 3496 13084 3505
rect 13136 3496 13138 3505
rect 13082 3431 13138 3440
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 800 12296 2246
rect 11978 96 12034 105
rect 11978 31 12034 40
rect 12254 0 12310 800
<< via2 >>
rect 1490 16360 1546 16416
rect 3072 14714 3128 14716
rect 3152 14714 3208 14716
rect 3232 14714 3288 14716
rect 3312 14714 3368 14716
rect 3072 14662 3118 14714
rect 3118 14662 3128 14714
rect 3152 14662 3182 14714
rect 3182 14662 3194 14714
rect 3194 14662 3208 14714
rect 3232 14662 3246 14714
rect 3246 14662 3258 14714
rect 3258 14662 3288 14714
rect 3312 14662 3322 14714
rect 3322 14662 3368 14714
rect 3072 14660 3128 14662
rect 3152 14660 3208 14662
rect 3232 14660 3288 14662
rect 3312 14660 3368 14662
rect 7304 14714 7360 14716
rect 7384 14714 7440 14716
rect 7464 14714 7520 14716
rect 7544 14714 7600 14716
rect 7304 14662 7350 14714
rect 7350 14662 7360 14714
rect 7384 14662 7414 14714
rect 7414 14662 7426 14714
rect 7426 14662 7440 14714
rect 7464 14662 7478 14714
rect 7478 14662 7490 14714
rect 7490 14662 7520 14714
rect 7544 14662 7554 14714
rect 7554 14662 7600 14714
rect 7304 14660 7360 14662
rect 7384 14660 7440 14662
rect 7464 14660 7520 14662
rect 7544 14660 7600 14662
rect 11536 14714 11592 14716
rect 11616 14714 11672 14716
rect 11696 14714 11752 14716
rect 11776 14714 11832 14716
rect 11536 14662 11582 14714
rect 11582 14662 11592 14714
rect 11616 14662 11646 14714
rect 11646 14662 11658 14714
rect 11658 14662 11672 14714
rect 11696 14662 11710 14714
rect 11710 14662 11722 14714
rect 11722 14662 11752 14714
rect 11776 14662 11786 14714
rect 11786 14662 11832 14714
rect 11536 14660 11592 14662
rect 11616 14660 11672 14662
rect 11696 14660 11752 14662
rect 11776 14660 11832 14662
rect 3072 13626 3128 13628
rect 3152 13626 3208 13628
rect 3232 13626 3288 13628
rect 3312 13626 3368 13628
rect 3072 13574 3118 13626
rect 3118 13574 3128 13626
rect 3152 13574 3182 13626
rect 3182 13574 3194 13626
rect 3194 13574 3208 13626
rect 3232 13574 3246 13626
rect 3246 13574 3258 13626
rect 3258 13574 3288 13626
rect 3312 13574 3322 13626
rect 3322 13574 3368 13626
rect 3072 13572 3128 13574
rect 3152 13572 3208 13574
rect 3232 13572 3288 13574
rect 3312 13572 3368 13574
rect 1490 12960 1546 13016
rect 3072 12538 3128 12540
rect 3152 12538 3208 12540
rect 3232 12538 3288 12540
rect 3312 12538 3368 12540
rect 3072 12486 3118 12538
rect 3118 12486 3128 12538
rect 3152 12486 3182 12538
rect 3182 12486 3194 12538
rect 3194 12486 3208 12538
rect 3232 12486 3246 12538
rect 3246 12486 3258 12538
rect 3258 12486 3288 12538
rect 3312 12486 3322 12538
rect 3322 12486 3368 12538
rect 3072 12484 3128 12486
rect 3152 12484 3208 12486
rect 3232 12484 3288 12486
rect 3312 12484 3368 12486
rect 3072 11450 3128 11452
rect 3152 11450 3208 11452
rect 3232 11450 3288 11452
rect 3312 11450 3368 11452
rect 3072 11398 3118 11450
rect 3118 11398 3128 11450
rect 3152 11398 3182 11450
rect 3182 11398 3194 11450
rect 3194 11398 3208 11450
rect 3232 11398 3246 11450
rect 3246 11398 3258 11450
rect 3258 11398 3288 11450
rect 3312 11398 3322 11450
rect 3322 11398 3368 11450
rect 3072 11396 3128 11398
rect 3152 11396 3208 11398
rect 3232 11396 3288 11398
rect 3312 11396 3368 11398
rect 5188 14170 5244 14172
rect 5268 14170 5324 14172
rect 5348 14170 5404 14172
rect 5428 14170 5484 14172
rect 5188 14118 5234 14170
rect 5234 14118 5244 14170
rect 5268 14118 5298 14170
rect 5298 14118 5310 14170
rect 5310 14118 5324 14170
rect 5348 14118 5362 14170
rect 5362 14118 5374 14170
rect 5374 14118 5404 14170
rect 5428 14118 5438 14170
rect 5438 14118 5484 14170
rect 5188 14116 5244 14118
rect 5268 14116 5324 14118
rect 5348 14116 5404 14118
rect 5428 14116 5484 14118
rect 5188 13082 5244 13084
rect 5268 13082 5324 13084
rect 5348 13082 5404 13084
rect 5428 13082 5484 13084
rect 5188 13030 5234 13082
rect 5234 13030 5244 13082
rect 5268 13030 5298 13082
rect 5298 13030 5310 13082
rect 5310 13030 5324 13082
rect 5348 13030 5362 13082
rect 5362 13030 5374 13082
rect 5374 13030 5404 13082
rect 5428 13030 5438 13082
rect 5438 13030 5484 13082
rect 5188 13028 5244 13030
rect 5268 13028 5324 13030
rect 5348 13028 5404 13030
rect 5428 13028 5484 13030
rect 5188 11994 5244 11996
rect 5268 11994 5324 11996
rect 5348 11994 5404 11996
rect 5428 11994 5484 11996
rect 5188 11942 5234 11994
rect 5234 11942 5244 11994
rect 5268 11942 5298 11994
rect 5298 11942 5310 11994
rect 5310 11942 5324 11994
rect 5348 11942 5362 11994
rect 5362 11942 5374 11994
rect 5374 11942 5404 11994
rect 5428 11942 5438 11994
rect 5438 11942 5484 11994
rect 5188 11940 5244 11942
rect 5268 11940 5324 11942
rect 5348 11940 5404 11942
rect 5428 11940 5484 11942
rect 1398 9560 1454 9616
rect 1490 6160 1546 6216
rect 1490 2796 1492 2816
rect 1492 2796 1544 2816
rect 1544 2796 1546 2816
rect 1490 2760 1546 2796
rect 3072 10362 3128 10364
rect 3152 10362 3208 10364
rect 3232 10362 3288 10364
rect 3312 10362 3368 10364
rect 3072 10310 3118 10362
rect 3118 10310 3128 10362
rect 3152 10310 3182 10362
rect 3182 10310 3194 10362
rect 3194 10310 3208 10362
rect 3232 10310 3246 10362
rect 3246 10310 3258 10362
rect 3258 10310 3288 10362
rect 3312 10310 3322 10362
rect 3322 10310 3368 10362
rect 3072 10308 3128 10310
rect 3152 10308 3208 10310
rect 3232 10308 3288 10310
rect 3312 10308 3368 10310
rect 3072 9274 3128 9276
rect 3152 9274 3208 9276
rect 3232 9274 3288 9276
rect 3312 9274 3368 9276
rect 3072 9222 3118 9274
rect 3118 9222 3128 9274
rect 3152 9222 3182 9274
rect 3182 9222 3194 9274
rect 3194 9222 3208 9274
rect 3232 9222 3246 9274
rect 3246 9222 3258 9274
rect 3258 9222 3288 9274
rect 3312 9222 3322 9274
rect 3322 9222 3368 9274
rect 3072 9220 3128 9222
rect 3152 9220 3208 9222
rect 3232 9220 3288 9222
rect 3312 9220 3368 9222
rect 5188 10906 5244 10908
rect 5268 10906 5324 10908
rect 5348 10906 5404 10908
rect 5428 10906 5484 10908
rect 5188 10854 5234 10906
rect 5234 10854 5244 10906
rect 5268 10854 5298 10906
rect 5298 10854 5310 10906
rect 5310 10854 5324 10906
rect 5348 10854 5362 10906
rect 5362 10854 5374 10906
rect 5374 10854 5404 10906
rect 5428 10854 5438 10906
rect 5438 10854 5484 10906
rect 5188 10852 5244 10854
rect 5268 10852 5324 10854
rect 5348 10852 5404 10854
rect 5428 10852 5484 10854
rect 7304 13626 7360 13628
rect 7384 13626 7440 13628
rect 7464 13626 7520 13628
rect 7544 13626 7600 13628
rect 7304 13574 7350 13626
rect 7350 13574 7360 13626
rect 7384 13574 7414 13626
rect 7414 13574 7426 13626
rect 7426 13574 7440 13626
rect 7464 13574 7478 13626
rect 7478 13574 7490 13626
rect 7490 13574 7520 13626
rect 7544 13574 7554 13626
rect 7554 13574 7600 13626
rect 7304 13572 7360 13574
rect 7384 13572 7440 13574
rect 7464 13572 7520 13574
rect 7544 13572 7600 13574
rect 3072 8186 3128 8188
rect 3152 8186 3208 8188
rect 3232 8186 3288 8188
rect 3312 8186 3368 8188
rect 3072 8134 3118 8186
rect 3118 8134 3128 8186
rect 3152 8134 3182 8186
rect 3182 8134 3194 8186
rect 3194 8134 3208 8186
rect 3232 8134 3246 8186
rect 3246 8134 3258 8186
rect 3258 8134 3288 8186
rect 3312 8134 3322 8186
rect 3322 8134 3368 8186
rect 3072 8132 3128 8134
rect 3152 8132 3208 8134
rect 3232 8132 3288 8134
rect 3312 8132 3368 8134
rect 3072 7098 3128 7100
rect 3152 7098 3208 7100
rect 3232 7098 3288 7100
rect 3312 7098 3368 7100
rect 3072 7046 3118 7098
rect 3118 7046 3128 7098
rect 3152 7046 3182 7098
rect 3182 7046 3194 7098
rect 3194 7046 3208 7098
rect 3232 7046 3246 7098
rect 3246 7046 3258 7098
rect 3258 7046 3288 7098
rect 3312 7046 3322 7098
rect 3322 7046 3368 7098
rect 3072 7044 3128 7046
rect 3152 7044 3208 7046
rect 3232 7044 3288 7046
rect 3312 7044 3368 7046
rect 5188 9818 5244 9820
rect 5268 9818 5324 9820
rect 5348 9818 5404 9820
rect 5428 9818 5484 9820
rect 5188 9766 5234 9818
rect 5234 9766 5244 9818
rect 5268 9766 5298 9818
rect 5298 9766 5310 9818
rect 5310 9766 5324 9818
rect 5348 9766 5362 9818
rect 5362 9766 5374 9818
rect 5374 9766 5404 9818
rect 5428 9766 5438 9818
rect 5438 9766 5484 9818
rect 5188 9764 5244 9766
rect 5268 9764 5324 9766
rect 5348 9764 5404 9766
rect 5428 9764 5484 9766
rect 7304 12538 7360 12540
rect 7384 12538 7440 12540
rect 7464 12538 7520 12540
rect 7544 12538 7600 12540
rect 7304 12486 7350 12538
rect 7350 12486 7360 12538
rect 7384 12486 7414 12538
rect 7414 12486 7426 12538
rect 7426 12486 7440 12538
rect 7464 12486 7478 12538
rect 7478 12486 7490 12538
rect 7490 12486 7520 12538
rect 7544 12486 7554 12538
rect 7554 12486 7600 12538
rect 7304 12484 7360 12486
rect 7384 12484 7440 12486
rect 7464 12484 7520 12486
rect 7544 12484 7600 12486
rect 7304 11450 7360 11452
rect 7384 11450 7440 11452
rect 7464 11450 7520 11452
rect 7544 11450 7600 11452
rect 7304 11398 7350 11450
rect 7350 11398 7360 11450
rect 7384 11398 7414 11450
rect 7414 11398 7426 11450
rect 7426 11398 7440 11450
rect 7464 11398 7478 11450
rect 7478 11398 7490 11450
rect 7490 11398 7520 11450
rect 7544 11398 7554 11450
rect 7554 11398 7600 11450
rect 7304 11396 7360 11398
rect 7384 11396 7440 11398
rect 7464 11396 7520 11398
rect 7544 11396 7600 11398
rect 5188 8730 5244 8732
rect 5268 8730 5324 8732
rect 5348 8730 5404 8732
rect 5428 8730 5484 8732
rect 5188 8678 5234 8730
rect 5234 8678 5244 8730
rect 5268 8678 5298 8730
rect 5298 8678 5310 8730
rect 5310 8678 5324 8730
rect 5348 8678 5362 8730
rect 5362 8678 5374 8730
rect 5374 8678 5404 8730
rect 5428 8678 5438 8730
rect 5438 8678 5484 8730
rect 5188 8676 5244 8678
rect 5268 8676 5324 8678
rect 5348 8676 5404 8678
rect 5428 8676 5484 8678
rect 3072 6010 3128 6012
rect 3152 6010 3208 6012
rect 3232 6010 3288 6012
rect 3312 6010 3368 6012
rect 3072 5958 3118 6010
rect 3118 5958 3128 6010
rect 3152 5958 3182 6010
rect 3182 5958 3194 6010
rect 3194 5958 3208 6010
rect 3232 5958 3246 6010
rect 3246 5958 3258 6010
rect 3258 5958 3288 6010
rect 3312 5958 3322 6010
rect 3322 5958 3368 6010
rect 3072 5956 3128 5958
rect 3152 5956 3208 5958
rect 3232 5956 3288 5958
rect 3312 5956 3368 5958
rect 3072 4922 3128 4924
rect 3152 4922 3208 4924
rect 3232 4922 3288 4924
rect 3312 4922 3368 4924
rect 3072 4870 3118 4922
rect 3118 4870 3128 4922
rect 3152 4870 3182 4922
rect 3182 4870 3194 4922
rect 3194 4870 3208 4922
rect 3232 4870 3246 4922
rect 3246 4870 3258 4922
rect 3258 4870 3288 4922
rect 3312 4870 3322 4922
rect 3322 4870 3368 4922
rect 3072 4868 3128 4870
rect 3152 4868 3208 4870
rect 3232 4868 3288 4870
rect 3312 4868 3368 4870
rect 5188 7642 5244 7644
rect 5268 7642 5324 7644
rect 5348 7642 5404 7644
rect 5428 7642 5484 7644
rect 5188 7590 5234 7642
rect 5234 7590 5244 7642
rect 5268 7590 5298 7642
rect 5298 7590 5310 7642
rect 5310 7590 5324 7642
rect 5348 7590 5362 7642
rect 5362 7590 5374 7642
rect 5374 7590 5404 7642
rect 5428 7590 5438 7642
rect 5438 7590 5484 7642
rect 5188 7588 5244 7590
rect 5268 7588 5324 7590
rect 5348 7588 5404 7590
rect 5428 7588 5484 7590
rect 5188 6554 5244 6556
rect 5268 6554 5324 6556
rect 5348 6554 5404 6556
rect 5428 6554 5484 6556
rect 5188 6502 5234 6554
rect 5234 6502 5244 6554
rect 5268 6502 5298 6554
rect 5298 6502 5310 6554
rect 5310 6502 5324 6554
rect 5348 6502 5362 6554
rect 5362 6502 5374 6554
rect 5374 6502 5404 6554
rect 5428 6502 5438 6554
rect 5438 6502 5484 6554
rect 5188 6500 5244 6502
rect 5268 6500 5324 6502
rect 5348 6500 5404 6502
rect 5428 6500 5484 6502
rect 7304 10362 7360 10364
rect 7384 10362 7440 10364
rect 7464 10362 7520 10364
rect 7544 10362 7600 10364
rect 7304 10310 7350 10362
rect 7350 10310 7360 10362
rect 7384 10310 7414 10362
rect 7414 10310 7426 10362
rect 7426 10310 7440 10362
rect 7464 10310 7478 10362
rect 7478 10310 7490 10362
rect 7490 10310 7520 10362
rect 7544 10310 7554 10362
rect 7554 10310 7600 10362
rect 7304 10308 7360 10310
rect 7384 10308 7440 10310
rect 7464 10308 7520 10310
rect 7544 10308 7600 10310
rect 7304 9274 7360 9276
rect 7384 9274 7440 9276
rect 7464 9274 7520 9276
rect 7544 9274 7600 9276
rect 7304 9222 7350 9274
rect 7350 9222 7360 9274
rect 7384 9222 7414 9274
rect 7414 9222 7426 9274
rect 7426 9222 7440 9274
rect 7464 9222 7478 9274
rect 7478 9222 7490 9274
rect 7490 9222 7520 9274
rect 7544 9222 7554 9274
rect 7554 9222 7600 9274
rect 7304 9220 7360 9222
rect 7384 9220 7440 9222
rect 7464 9220 7520 9222
rect 7544 9220 7600 9222
rect 7304 8186 7360 8188
rect 7384 8186 7440 8188
rect 7464 8186 7520 8188
rect 7544 8186 7600 8188
rect 7304 8134 7350 8186
rect 7350 8134 7360 8186
rect 7384 8134 7414 8186
rect 7414 8134 7426 8186
rect 7426 8134 7440 8186
rect 7464 8134 7478 8186
rect 7478 8134 7490 8186
rect 7490 8134 7520 8186
rect 7544 8134 7554 8186
rect 7554 8134 7600 8186
rect 7304 8132 7360 8134
rect 7384 8132 7440 8134
rect 7464 8132 7520 8134
rect 7544 8132 7600 8134
rect 7304 7098 7360 7100
rect 7384 7098 7440 7100
rect 7464 7098 7520 7100
rect 7544 7098 7600 7100
rect 7304 7046 7350 7098
rect 7350 7046 7360 7098
rect 7384 7046 7414 7098
rect 7414 7046 7426 7098
rect 7426 7046 7440 7098
rect 7464 7046 7478 7098
rect 7478 7046 7490 7098
rect 7490 7046 7520 7098
rect 7544 7046 7554 7098
rect 7554 7046 7600 7098
rect 7304 7044 7360 7046
rect 7384 7044 7440 7046
rect 7464 7044 7520 7046
rect 7544 7044 7600 7046
rect 5188 5466 5244 5468
rect 5268 5466 5324 5468
rect 5348 5466 5404 5468
rect 5428 5466 5484 5468
rect 5188 5414 5234 5466
rect 5234 5414 5244 5466
rect 5268 5414 5298 5466
rect 5298 5414 5310 5466
rect 5310 5414 5324 5466
rect 5348 5414 5362 5466
rect 5362 5414 5374 5466
rect 5374 5414 5404 5466
rect 5428 5414 5438 5466
rect 5438 5414 5484 5466
rect 5188 5412 5244 5414
rect 5268 5412 5324 5414
rect 5348 5412 5404 5414
rect 5428 5412 5484 5414
rect 5188 4378 5244 4380
rect 5268 4378 5324 4380
rect 5348 4378 5404 4380
rect 5428 4378 5484 4380
rect 5188 4326 5234 4378
rect 5234 4326 5244 4378
rect 5268 4326 5298 4378
rect 5298 4326 5310 4378
rect 5310 4326 5324 4378
rect 5348 4326 5362 4378
rect 5362 4326 5374 4378
rect 5374 4326 5404 4378
rect 5428 4326 5438 4378
rect 5438 4326 5484 4378
rect 5188 4324 5244 4326
rect 5268 4324 5324 4326
rect 5348 4324 5404 4326
rect 5428 4324 5484 4326
rect 3072 3834 3128 3836
rect 3152 3834 3208 3836
rect 3232 3834 3288 3836
rect 3312 3834 3368 3836
rect 3072 3782 3118 3834
rect 3118 3782 3128 3834
rect 3152 3782 3182 3834
rect 3182 3782 3194 3834
rect 3194 3782 3208 3834
rect 3232 3782 3246 3834
rect 3246 3782 3258 3834
rect 3258 3782 3288 3834
rect 3312 3782 3322 3834
rect 3322 3782 3368 3834
rect 3072 3780 3128 3782
rect 3152 3780 3208 3782
rect 3232 3780 3288 3782
rect 3312 3780 3368 3782
rect 5188 3290 5244 3292
rect 5268 3290 5324 3292
rect 5348 3290 5404 3292
rect 5428 3290 5484 3292
rect 5188 3238 5234 3290
rect 5234 3238 5244 3290
rect 5268 3238 5298 3290
rect 5298 3238 5310 3290
rect 5310 3238 5324 3290
rect 5348 3238 5362 3290
rect 5362 3238 5374 3290
rect 5374 3238 5404 3290
rect 5428 3238 5438 3290
rect 5438 3238 5484 3290
rect 5188 3236 5244 3238
rect 5268 3236 5324 3238
rect 5348 3236 5404 3238
rect 5428 3236 5484 3238
rect 3072 2746 3128 2748
rect 3152 2746 3208 2748
rect 3232 2746 3288 2748
rect 3312 2746 3368 2748
rect 3072 2694 3118 2746
rect 3118 2694 3128 2746
rect 3152 2694 3182 2746
rect 3182 2694 3194 2746
rect 3194 2694 3208 2746
rect 3232 2694 3246 2746
rect 3246 2694 3258 2746
rect 3258 2694 3288 2746
rect 3312 2694 3322 2746
rect 3322 2694 3368 2746
rect 3072 2692 3128 2694
rect 3152 2692 3208 2694
rect 3232 2692 3288 2694
rect 3312 2692 3368 2694
rect 7304 6010 7360 6012
rect 7384 6010 7440 6012
rect 7464 6010 7520 6012
rect 7544 6010 7600 6012
rect 7304 5958 7350 6010
rect 7350 5958 7360 6010
rect 7384 5958 7414 6010
rect 7414 5958 7426 6010
rect 7426 5958 7440 6010
rect 7464 5958 7478 6010
rect 7478 5958 7490 6010
rect 7490 5958 7520 6010
rect 7544 5958 7554 6010
rect 7554 5958 7600 6010
rect 7304 5956 7360 5958
rect 7384 5956 7440 5958
rect 7464 5956 7520 5958
rect 7544 5956 7600 5958
rect 9420 14170 9476 14172
rect 9500 14170 9556 14172
rect 9580 14170 9636 14172
rect 9660 14170 9716 14172
rect 9420 14118 9466 14170
rect 9466 14118 9476 14170
rect 9500 14118 9530 14170
rect 9530 14118 9542 14170
rect 9542 14118 9556 14170
rect 9580 14118 9594 14170
rect 9594 14118 9606 14170
rect 9606 14118 9636 14170
rect 9660 14118 9670 14170
rect 9670 14118 9716 14170
rect 9420 14116 9476 14118
rect 9500 14116 9556 14118
rect 9580 14116 9636 14118
rect 9660 14116 9716 14118
rect 9420 13082 9476 13084
rect 9500 13082 9556 13084
rect 9580 13082 9636 13084
rect 9660 13082 9716 13084
rect 9420 13030 9466 13082
rect 9466 13030 9476 13082
rect 9500 13030 9530 13082
rect 9530 13030 9542 13082
rect 9542 13030 9556 13082
rect 9580 13030 9594 13082
rect 9594 13030 9606 13082
rect 9606 13030 9636 13082
rect 9660 13030 9670 13082
rect 9670 13030 9716 13082
rect 9420 13028 9476 13030
rect 9500 13028 9556 13030
rect 9580 13028 9636 13030
rect 9660 13028 9716 13030
rect 9420 11994 9476 11996
rect 9500 11994 9556 11996
rect 9580 11994 9636 11996
rect 9660 11994 9716 11996
rect 9420 11942 9466 11994
rect 9466 11942 9476 11994
rect 9500 11942 9530 11994
rect 9530 11942 9542 11994
rect 9542 11942 9556 11994
rect 9580 11942 9594 11994
rect 9594 11942 9606 11994
rect 9606 11942 9636 11994
rect 9660 11942 9670 11994
rect 9670 11942 9716 11994
rect 9420 11940 9476 11942
rect 9500 11940 9556 11942
rect 9580 11940 9636 11942
rect 9660 11940 9716 11942
rect 9420 10906 9476 10908
rect 9500 10906 9556 10908
rect 9580 10906 9636 10908
rect 9660 10906 9716 10908
rect 9420 10854 9466 10906
rect 9466 10854 9476 10906
rect 9500 10854 9530 10906
rect 9530 10854 9542 10906
rect 9542 10854 9556 10906
rect 9580 10854 9594 10906
rect 9594 10854 9606 10906
rect 9606 10854 9636 10906
rect 9660 10854 9670 10906
rect 9670 10854 9716 10906
rect 9420 10852 9476 10854
rect 9500 10852 9556 10854
rect 9580 10852 9636 10854
rect 9660 10852 9716 10854
rect 11536 13626 11592 13628
rect 11616 13626 11672 13628
rect 11696 13626 11752 13628
rect 11776 13626 11832 13628
rect 11536 13574 11582 13626
rect 11582 13574 11592 13626
rect 11616 13574 11646 13626
rect 11646 13574 11658 13626
rect 11658 13574 11672 13626
rect 11696 13574 11710 13626
rect 11710 13574 11722 13626
rect 11722 13574 11752 13626
rect 11776 13574 11786 13626
rect 11786 13574 11832 13626
rect 11536 13572 11592 13574
rect 11616 13572 11672 13574
rect 11696 13572 11752 13574
rect 11776 13572 11832 13574
rect 11536 12538 11592 12540
rect 11616 12538 11672 12540
rect 11696 12538 11752 12540
rect 11776 12538 11832 12540
rect 11536 12486 11582 12538
rect 11582 12486 11592 12538
rect 11616 12486 11646 12538
rect 11646 12486 11658 12538
rect 11658 12486 11672 12538
rect 11696 12486 11710 12538
rect 11710 12486 11722 12538
rect 11722 12486 11752 12538
rect 11776 12486 11786 12538
rect 11786 12486 11832 12538
rect 11536 12484 11592 12486
rect 11616 12484 11672 12486
rect 11696 12484 11752 12486
rect 11776 12484 11832 12486
rect 11536 11450 11592 11452
rect 11616 11450 11672 11452
rect 11696 11450 11752 11452
rect 11776 11450 11832 11452
rect 11536 11398 11582 11450
rect 11582 11398 11592 11450
rect 11616 11398 11646 11450
rect 11646 11398 11658 11450
rect 11658 11398 11672 11450
rect 11696 11398 11710 11450
rect 11710 11398 11722 11450
rect 11722 11398 11752 11450
rect 11776 11398 11786 11450
rect 11786 11398 11832 11450
rect 11536 11396 11592 11398
rect 11616 11396 11672 11398
rect 11696 11396 11752 11398
rect 11776 11396 11832 11398
rect 9420 9818 9476 9820
rect 9500 9818 9556 9820
rect 9580 9818 9636 9820
rect 9660 9818 9716 9820
rect 9420 9766 9466 9818
rect 9466 9766 9476 9818
rect 9500 9766 9530 9818
rect 9530 9766 9542 9818
rect 9542 9766 9556 9818
rect 9580 9766 9594 9818
rect 9594 9766 9606 9818
rect 9606 9766 9636 9818
rect 9660 9766 9670 9818
rect 9670 9766 9716 9818
rect 9420 9764 9476 9766
rect 9500 9764 9556 9766
rect 9580 9764 9636 9766
rect 9660 9764 9716 9766
rect 11536 10362 11592 10364
rect 11616 10362 11672 10364
rect 11696 10362 11752 10364
rect 11776 10362 11832 10364
rect 11536 10310 11582 10362
rect 11582 10310 11592 10362
rect 11616 10310 11646 10362
rect 11646 10310 11658 10362
rect 11658 10310 11672 10362
rect 11696 10310 11710 10362
rect 11710 10310 11722 10362
rect 11722 10310 11752 10362
rect 11776 10310 11786 10362
rect 11786 10310 11832 10362
rect 11536 10308 11592 10310
rect 11616 10308 11672 10310
rect 11696 10308 11752 10310
rect 11776 10308 11832 10310
rect 11536 9274 11592 9276
rect 11616 9274 11672 9276
rect 11696 9274 11752 9276
rect 11776 9274 11832 9276
rect 11536 9222 11582 9274
rect 11582 9222 11592 9274
rect 11616 9222 11646 9274
rect 11646 9222 11658 9274
rect 11658 9222 11672 9274
rect 11696 9222 11710 9274
rect 11710 9222 11722 9274
rect 11722 9222 11752 9274
rect 11776 9222 11786 9274
rect 11786 9222 11832 9274
rect 11536 9220 11592 9222
rect 11616 9220 11672 9222
rect 11696 9220 11752 9222
rect 11776 9220 11832 9222
rect 9420 8730 9476 8732
rect 9500 8730 9556 8732
rect 9580 8730 9636 8732
rect 9660 8730 9716 8732
rect 9420 8678 9466 8730
rect 9466 8678 9476 8730
rect 9500 8678 9530 8730
rect 9530 8678 9542 8730
rect 9542 8678 9556 8730
rect 9580 8678 9594 8730
rect 9594 8678 9606 8730
rect 9606 8678 9636 8730
rect 9660 8678 9670 8730
rect 9670 8678 9716 8730
rect 9420 8676 9476 8678
rect 9500 8676 9556 8678
rect 9580 8676 9636 8678
rect 9660 8676 9716 8678
rect 11536 8186 11592 8188
rect 11616 8186 11672 8188
rect 11696 8186 11752 8188
rect 11776 8186 11832 8188
rect 11536 8134 11582 8186
rect 11582 8134 11592 8186
rect 11616 8134 11646 8186
rect 11646 8134 11658 8186
rect 11658 8134 11672 8186
rect 11696 8134 11710 8186
rect 11710 8134 11722 8186
rect 11722 8134 11752 8186
rect 11776 8134 11786 8186
rect 11786 8134 11832 8186
rect 11536 8132 11592 8134
rect 11616 8132 11672 8134
rect 11696 8132 11752 8134
rect 11776 8132 11832 8134
rect 12990 13676 12992 13696
rect 12992 13676 13044 13696
rect 13044 13676 13046 13696
rect 12990 13640 13046 13676
rect 9420 7642 9476 7644
rect 9500 7642 9556 7644
rect 9580 7642 9636 7644
rect 9660 7642 9716 7644
rect 9420 7590 9466 7642
rect 9466 7590 9476 7642
rect 9500 7590 9530 7642
rect 9530 7590 9542 7642
rect 9542 7590 9556 7642
rect 9580 7590 9594 7642
rect 9594 7590 9606 7642
rect 9606 7590 9636 7642
rect 9660 7590 9670 7642
rect 9670 7590 9716 7642
rect 9420 7588 9476 7590
rect 9500 7588 9556 7590
rect 9580 7588 9636 7590
rect 9660 7588 9716 7590
rect 11536 7098 11592 7100
rect 11616 7098 11672 7100
rect 11696 7098 11752 7100
rect 11776 7098 11832 7100
rect 11536 7046 11582 7098
rect 11582 7046 11592 7098
rect 11616 7046 11646 7098
rect 11646 7046 11658 7098
rect 11658 7046 11672 7098
rect 11696 7046 11710 7098
rect 11710 7046 11722 7098
rect 11722 7046 11752 7098
rect 11776 7046 11786 7098
rect 11786 7046 11832 7098
rect 11536 7044 11592 7046
rect 11616 7044 11672 7046
rect 11696 7044 11752 7046
rect 11776 7044 11832 7046
rect 9420 6554 9476 6556
rect 9500 6554 9556 6556
rect 9580 6554 9636 6556
rect 9660 6554 9716 6556
rect 9420 6502 9466 6554
rect 9466 6502 9476 6554
rect 9500 6502 9530 6554
rect 9530 6502 9542 6554
rect 9542 6502 9556 6554
rect 9580 6502 9594 6554
rect 9594 6502 9606 6554
rect 9606 6502 9636 6554
rect 9660 6502 9670 6554
rect 9670 6502 9716 6554
rect 9420 6500 9476 6502
rect 9500 6500 9556 6502
rect 9580 6500 9636 6502
rect 9660 6500 9716 6502
rect 11536 6010 11592 6012
rect 11616 6010 11672 6012
rect 11696 6010 11752 6012
rect 11776 6010 11832 6012
rect 11536 5958 11582 6010
rect 11582 5958 11592 6010
rect 11616 5958 11646 6010
rect 11646 5958 11658 6010
rect 11658 5958 11672 6010
rect 11696 5958 11710 6010
rect 11710 5958 11722 6010
rect 11722 5958 11752 6010
rect 11776 5958 11786 6010
rect 11786 5958 11832 6010
rect 11536 5956 11592 5958
rect 11616 5956 11672 5958
rect 11696 5956 11752 5958
rect 11776 5956 11832 5958
rect 7304 4922 7360 4924
rect 7384 4922 7440 4924
rect 7464 4922 7520 4924
rect 7544 4922 7600 4924
rect 7304 4870 7350 4922
rect 7350 4870 7360 4922
rect 7384 4870 7414 4922
rect 7414 4870 7426 4922
rect 7426 4870 7440 4922
rect 7464 4870 7478 4922
rect 7478 4870 7490 4922
rect 7490 4870 7520 4922
rect 7544 4870 7554 4922
rect 7554 4870 7600 4922
rect 7304 4868 7360 4870
rect 7384 4868 7440 4870
rect 7464 4868 7520 4870
rect 7544 4868 7600 4870
rect 7304 3834 7360 3836
rect 7384 3834 7440 3836
rect 7464 3834 7520 3836
rect 7544 3834 7600 3836
rect 7304 3782 7350 3834
rect 7350 3782 7360 3834
rect 7384 3782 7414 3834
rect 7414 3782 7426 3834
rect 7426 3782 7440 3834
rect 7464 3782 7478 3834
rect 7478 3782 7490 3834
rect 7490 3782 7520 3834
rect 7544 3782 7554 3834
rect 7554 3782 7600 3834
rect 7304 3780 7360 3782
rect 7384 3780 7440 3782
rect 7464 3780 7520 3782
rect 7544 3780 7600 3782
rect 7304 2746 7360 2748
rect 7384 2746 7440 2748
rect 7464 2746 7520 2748
rect 7544 2746 7600 2748
rect 7304 2694 7350 2746
rect 7350 2694 7360 2746
rect 7384 2694 7414 2746
rect 7414 2694 7426 2746
rect 7426 2694 7440 2746
rect 7464 2694 7478 2746
rect 7478 2694 7490 2746
rect 7490 2694 7520 2746
rect 7544 2694 7554 2746
rect 7554 2694 7600 2746
rect 7304 2692 7360 2694
rect 7384 2692 7440 2694
rect 7464 2692 7520 2694
rect 7544 2692 7600 2694
rect 9420 5466 9476 5468
rect 9500 5466 9556 5468
rect 9580 5466 9636 5468
rect 9660 5466 9716 5468
rect 9420 5414 9466 5466
rect 9466 5414 9476 5466
rect 9500 5414 9530 5466
rect 9530 5414 9542 5466
rect 9542 5414 9556 5466
rect 9580 5414 9594 5466
rect 9594 5414 9606 5466
rect 9606 5414 9636 5466
rect 9660 5414 9670 5466
rect 9670 5414 9716 5466
rect 9420 5412 9476 5414
rect 9500 5412 9556 5414
rect 9580 5412 9636 5414
rect 9660 5412 9716 5414
rect 11536 4922 11592 4924
rect 11616 4922 11672 4924
rect 11696 4922 11752 4924
rect 11776 4922 11832 4924
rect 11536 4870 11582 4922
rect 11582 4870 11592 4922
rect 11616 4870 11646 4922
rect 11646 4870 11658 4922
rect 11658 4870 11672 4922
rect 11696 4870 11710 4922
rect 11710 4870 11722 4922
rect 11722 4870 11752 4922
rect 11776 4870 11786 4922
rect 11786 4870 11832 4922
rect 11536 4868 11592 4870
rect 11616 4868 11672 4870
rect 11696 4868 11752 4870
rect 11776 4868 11832 4870
rect 9420 4378 9476 4380
rect 9500 4378 9556 4380
rect 9580 4378 9636 4380
rect 9660 4378 9716 4380
rect 9420 4326 9466 4378
rect 9466 4326 9476 4378
rect 9500 4326 9530 4378
rect 9530 4326 9542 4378
rect 9542 4326 9556 4378
rect 9580 4326 9594 4378
rect 9594 4326 9606 4378
rect 9606 4326 9636 4378
rect 9660 4326 9670 4378
rect 9670 4326 9716 4378
rect 9420 4324 9476 4326
rect 9500 4324 9556 4326
rect 9580 4324 9636 4326
rect 9660 4324 9716 4326
rect 11536 3834 11592 3836
rect 11616 3834 11672 3836
rect 11696 3834 11752 3836
rect 11776 3834 11832 3836
rect 11536 3782 11582 3834
rect 11582 3782 11592 3834
rect 11616 3782 11646 3834
rect 11646 3782 11658 3834
rect 11658 3782 11672 3834
rect 11696 3782 11710 3834
rect 11710 3782 11722 3834
rect 11722 3782 11752 3834
rect 11776 3782 11786 3834
rect 11786 3782 11832 3834
rect 11536 3780 11592 3782
rect 11616 3780 11672 3782
rect 11696 3780 11752 3782
rect 11776 3780 11832 3782
rect 9420 3290 9476 3292
rect 9500 3290 9556 3292
rect 9580 3290 9636 3292
rect 9660 3290 9716 3292
rect 9420 3238 9466 3290
rect 9466 3238 9476 3290
rect 9500 3238 9530 3290
rect 9530 3238 9542 3290
rect 9542 3238 9556 3290
rect 9580 3238 9594 3290
rect 9594 3238 9606 3290
rect 9606 3238 9636 3290
rect 9660 3238 9670 3290
rect 9670 3238 9716 3290
rect 9420 3236 9476 3238
rect 9500 3236 9556 3238
rect 9580 3236 9636 3238
rect 9660 3236 9716 3238
rect 11536 2746 11592 2748
rect 11616 2746 11672 2748
rect 11696 2746 11752 2748
rect 11776 2746 11832 2748
rect 11536 2694 11582 2746
rect 11582 2694 11592 2746
rect 11616 2694 11646 2746
rect 11646 2694 11658 2746
rect 11658 2694 11672 2746
rect 11696 2694 11710 2746
rect 11710 2694 11722 2746
rect 11722 2694 11752 2746
rect 11776 2694 11786 2746
rect 11786 2694 11832 2746
rect 11536 2692 11592 2694
rect 11616 2692 11672 2694
rect 11696 2692 11752 2694
rect 11776 2692 11832 2694
rect 5188 2202 5244 2204
rect 5268 2202 5324 2204
rect 5348 2202 5404 2204
rect 5428 2202 5484 2204
rect 5188 2150 5234 2202
rect 5234 2150 5244 2202
rect 5268 2150 5298 2202
rect 5298 2150 5310 2202
rect 5310 2150 5324 2202
rect 5348 2150 5362 2202
rect 5362 2150 5374 2202
rect 5374 2150 5404 2202
rect 5428 2150 5438 2202
rect 5438 2150 5484 2202
rect 5188 2148 5244 2150
rect 5268 2148 5324 2150
rect 5348 2148 5404 2150
rect 5428 2148 5484 2150
rect 9420 2202 9476 2204
rect 9500 2202 9556 2204
rect 9580 2202 9636 2204
rect 9660 2202 9716 2204
rect 9420 2150 9466 2202
rect 9466 2150 9476 2202
rect 9500 2150 9530 2202
rect 9530 2150 9542 2202
rect 9542 2150 9556 2202
rect 9580 2150 9594 2202
rect 9594 2150 9606 2202
rect 9606 2150 9636 2202
rect 9660 2150 9670 2202
rect 9670 2150 9716 2202
rect 9420 2148 9476 2150
rect 9500 2148 9556 2150
rect 9580 2148 9636 2150
rect 9660 2148 9716 2150
rect 12990 10240 13046 10296
rect 13082 6840 13138 6896
rect 13082 3476 13084 3496
rect 13084 3476 13136 3496
rect 13136 3476 13138 3496
rect 13082 3440 13138 3476
rect 11978 40 12034 96
<< metal3 >>
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 3060 14720 3380 14721
rect 3060 14656 3068 14720
rect 3132 14656 3148 14720
rect 3212 14656 3228 14720
rect 3292 14656 3308 14720
rect 3372 14656 3380 14720
rect 3060 14655 3380 14656
rect 7292 14720 7612 14721
rect 7292 14656 7300 14720
rect 7364 14656 7380 14720
rect 7444 14656 7460 14720
rect 7524 14656 7540 14720
rect 7604 14656 7612 14720
rect 7292 14655 7612 14656
rect 11524 14720 11844 14721
rect 11524 14656 11532 14720
rect 11596 14656 11612 14720
rect 11676 14656 11692 14720
rect 11756 14656 11772 14720
rect 11836 14656 11844 14720
rect 11524 14655 11844 14656
rect 5176 14176 5496 14177
rect 5176 14112 5184 14176
rect 5248 14112 5264 14176
rect 5328 14112 5344 14176
rect 5408 14112 5424 14176
rect 5488 14112 5496 14176
rect 5176 14111 5496 14112
rect 9408 14176 9728 14177
rect 9408 14112 9416 14176
rect 9480 14112 9496 14176
rect 9560 14112 9576 14176
rect 9640 14112 9656 14176
rect 9720 14112 9728 14176
rect 9408 14111 9728 14112
rect 12985 13698 13051 13701
rect 14181 13698 14981 13728
rect 12985 13696 14981 13698
rect 12985 13640 12990 13696
rect 13046 13640 14981 13696
rect 12985 13638 14981 13640
rect 12985 13635 13051 13638
rect 3060 13632 3380 13633
rect 3060 13568 3068 13632
rect 3132 13568 3148 13632
rect 3212 13568 3228 13632
rect 3292 13568 3308 13632
rect 3372 13568 3380 13632
rect 3060 13567 3380 13568
rect 7292 13632 7612 13633
rect 7292 13568 7300 13632
rect 7364 13568 7380 13632
rect 7444 13568 7460 13632
rect 7524 13568 7540 13632
rect 7604 13568 7612 13632
rect 7292 13567 7612 13568
rect 11524 13632 11844 13633
rect 11524 13568 11532 13632
rect 11596 13568 11612 13632
rect 11676 13568 11692 13632
rect 11756 13568 11772 13632
rect 11836 13568 11844 13632
rect 14181 13608 14981 13638
rect 11524 13567 11844 13568
rect 5176 13088 5496 13089
rect 0 13018 800 13048
rect 5176 13024 5184 13088
rect 5248 13024 5264 13088
rect 5328 13024 5344 13088
rect 5408 13024 5424 13088
rect 5488 13024 5496 13088
rect 5176 13023 5496 13024
rect 9408 13088 9728 13089
rect 9408 13024 9416 13088
rect 9480 13024 9496 13088
rect 9560 13024 9576 13088
rect 9640 13024 9656 13088
rect 9720 13024 9728 13088
rect 9408 13023 9728 13024
rect 1485 13018 1551 13021
rect 0 13016 1551 13018
rect 0 12960 1490 13016
rect 1546 12960 1551 13016
rect 0 12958 1551 12960
rect 0 12928 800 12958
rect 1485 12955 1551 12958
rect 3060 12544 3380 12545
rect 3060 12480 3068 12544
rect 3132 12480 3148 12544
rect 3212 12480 3228 12544
rect 3292 12480 3308 12544
rect 3372 12480 3380 12544
rect 3060 12479 3380 12480
rect 7292 12544 7612 12545
rect 7292 12480 7300 12544
rect 7364 12480 7380 12544
rect 7444 12480 7460 12544
rect 7524 12480 7540 12544
rect 7604 12480 7612 12544
rect 7292 12479 7612 12480
rect 11524 12544 11844 12545
rect 11524 12480 11532 12544
rect 11596 12480 11612 12544
rect 11676 12480 11692 12544
rect 11756 12480 11772 12544
rect 11836 12480 11844 12544
rect 11524 12479 11844 12480
rect 5176 12000 5496 12001
rect 5176 11936 5184 12000
rect 5248 11936 5264 12000
rect 5328 11936 5344 12000
rect 5408 11936 5424 12000
rect 5488 11936 5496 12000
rect 5176 11935 5496 11936
rect 9408 12000 9728 12001
rect 9408 11936 9416 12000
rect 9480 11936 9496 12000
rect 9560 11936 9576 12000
rect 9640 11936 9656 12000
rect 9720 11936 9728 12000
rect 9408 11935 9728 11936
rect 3060 11456 3380 11457
rect 3060 11392 3068 11456
rect 3132 11392 3148 11456
rect 3212 11392 3228 11456
rect 3292 11392 3308 11456
rect 3372 11392 3380 11456
rect 3060 11391 3380 11392
rect 7292 11456 7612 11457
rect 7292 11392 7300 11456
rect 7364 11392 7380 11456
rect 7444 11392 7460 11456
rect 7524 11392 7540 11456
rect 7604 11392 7612 11456
rect 7292 11391 7612 11392
rect 11524 11456 11844 11457
rect 11524 11392 11532 11456
rect 11596 11392 11612 11456
rect 11676 11392 11692 11456
rect 11756 11392 11772 11456
rect 11836 11392 11844 11456
rect 11524 11391 11844 11392
rect 5176 10912 5496 10913
rect 5176 10848 5184 10912
rect 5248 10848 5264 10912
rect 5328 10848 5344 10912
rect 5408 10848 5424 10912
rect 5488 10848 5496 10912
rect 5176 10847 5496 10848
rect 9408 10912 9728 10913
rect 9408 10848 9416 10912
rect 9480 10848 9496 10912
rect 9560 10848 9576 10912
rect 9640 10848 9656 10912
rect 9720 10848 9728 10912
rect 9408 10847 9728 10848
rect 3060 10368 3380 10369
rect 3060 10304 3068 10368
rect 3132 10304 3148 10368
rect 3212 10304 3228 10368
rect 3292 10304 3308 10368
rect 3372 10304 3380 10368
rect 3060 10303 3380 10304
rect 7292 10368 7612 10369
rect 7292 10304 7300 10368
rect 7364 10304 7380 10368
rect 7444 10304 7460 10368
rect 7524 10304 7540 10368
rect 7604 10304 7612 10368
rect 7292 10303 7612 10304
rect 11524 10368 11844 10369
rect 11524 10304 11532 10368
rect 11596 10304 11612 10368
rect 11676 10304 11692 10368
rect 11756 10304 11772 10368
rect 11836 10304 11844 10368
rect 11524 10303 11844 10304
rect 12985 10298 13051 10301
rect 14181 10298 14981 10328
rect 12985 10296 14981 10298
rect 12985 10240 12990 10296
rect 13046 10240 14981 10296
rect 12985 10238 14981 10240
rect 12985 10235 13051 10238
rect 14181 10208 14981 10238
rect 5176 9824 5496 9825
rect 5176 9760 5184 9824
rect 5248 9760 5264 9824
rect 5328 9760 5344 9824
rect 5408 9760 5424 9824
rect 5488 9760 5496 9824
rect 5176 9759 5496 9760
rect 9408 9824 9728 9825
rect 9408 9760 9416 9824
rect 9480 9760 9496 9824
rect 9560 9760 9576 9824
rect 9640 9760 9656 9824
rect 9720 9760 9728 9824
rect 9408 9759 9728 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 3060 9280 3380 9281
rect 3060 9216 3068 9280
rect 3132 9216 3148 9280
rect 3212 9216 3228 9280
rect 3292 9216 3308 9280
rect 3372 9216 3380 9280
rect 3060 9215 3380 9216
rect 7292 9280 7612 9281
rect 7292 9216 7300 9280
rect 7364 9216 7380 9280
rect 7444 9216 7460 9280
rect 7524 9216 7540 9280
rect 7604 9216 7612 9280
rect 7292 9215 7612 9216
rect 11524 9280 11844 9281
rect 11524 9216 11532 9280
rect 11596 9216 11612 9280
rect 11676 9216 11692 9280
rect 11756 9216 11772 9280
rect 11836 9216 11844 9280
rect 11524 9215 11844 9216
rect 5176 8736 5496 8737
rect 5176 8672 5184 8736
rect 5248 8672 5264 8736
rect 5328 8672 5344 8736
rect 5408 8672 5424 8736
rect 5488 8672 5496 8736
rect 5176 8671 5496 8672
rect 9408 8736 9728 8737
rect 9408 8672 9416 8736
rect 9480 8672 9496 8736
rect 9560 8672 9576 8736
rect 9640 8672 9656 8736
rect 9720 8672 9728 8736
rect 9408 8671 9728 8672
rect 3060 8192 3380 8193
rect 3060 8128 3068 8192
rect 3132 8128 3148 8192
rect 3212 8128 3228 8192
rect 3292 8128 3308 8192
rect 3372 8128 3380 8192
rect 3060 8127 3380 8128
rect 7292 8192 7612 8193
rect 7292 8128 7300 8192
rect 7364 8128 7380 8192
rect 7444 8128 7460 8192
rect 7524 8128 7540 8192
rect 7604 8128 7612 8192
rect 7292 8127 7612 8128
rect 11524 8192 11844 8193
rect 11524 8128 11532 8192
rect 11596 8128 11612 8192
rect 11676 8128 11692 8192
rect 11756 8128 11772 8192
rect 11836 8128 11844 8192
rect 11524 8127 11844 8128
rect 5176 7648 5496 7649
rect 5176 7584 5184 7648
rect 5248 7584 5264 7648
rect 5328 7584 5344 7648
rect 5408 7584 5424 7648
rect 5488 7584 5496 7648
rect 5176 7583 5496 7584
rect 9408 7648 9728 7649
rect 9408 7584 9416 7648
rect 9480 7584 9496 7648
rect 9560 7584 9576 7648
rect 9640 7584 9656 7648
rect 9720 7584 9728 7648
rect 9408 7583 9728 7584
rect 3060 7104 3380 7105
rect 3060 7040 3068 7104
rect 3132 7040 3148 7104
rect 3212 7040 3228 7104
rect 3292 7040 3308 7104
rect 3372 7040 3380 7104
rect 3060 7039 3380 7040
rect 7292 7104 7612 7105
rect 7292 7040 7300 7104
rect 7364 7040 7380 7104
rect 7444 7040 7460 7104
rect 7524 7040 7540 7104
rect 7604 7040 7612 7104
rect 7292 7039 7612 7040
rect 11524 7104 11844 7105
rect 11524 7040 11532 7104
rect 11596 7040 11612 7104
rect 11676 7040 11692 7104
rect 11756 7040 11772 7104
rect 11836 7040 11844 7104
rect 11524 7039 11844 7040
rect 13077 6898 13143 6901
rect 14181 6898 14981 6928
rect 13077 6896 14981 6898
rect 13077 6840 13082 6896
rect 13138 6840 14981 6896
rect 13077 6838 14981 6840
rect 13077 6835 13143 6838
rect 14181 6808 14981 6838
rect 5176 6560 5496 6561
rect 5176 6496 5184 6560
rect 5248 6496 5264 6560
rect 5328 6496 5344 6560
rect 5408 6496 5424 6560
rect 5488 6496 5496 6560
rect 5176 6495 5496 6496
rect 9408 6560 9728 6561
rect 9408 6496 9416 6560
rect 9480 6496 9496 6560
rect 9560 6496 9576 6560
rect 9640 6496 9656 6560
rect 9720 6496 9728 6560
rect 9408 6495 9728 6496
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 3060 6016 3380 6017
rect 3060 5952 3068 6016
rect 3132 5952 3148 6016
rect 3212 5952 3228 6016
rect 3292 5952 3308 6016
rect 3372 5952 3380 6016
rect 3060 5951 3380 5952
rect 7292 6016 7612 6017
rect 7292 5952 7300 6016
rect 7364 5952 7380 6016
rect 7444 5952 7460 6016
rect 7524 5952 7540 6016
rect 7604 5952 7612 6016
rect 7292 5951 7612 5952
rect 11524 6016 11844 6017
rect 11524 5952 11532 6016
rect 11596 5952 11612 6016
rect 11676 5952 11692 6016
rect 11756 5952 11772 6016
rect 11836 5952 11844 6016
rect 11524 5951 11844 5952
rect 5176 5472 5496 5473
rect 5176 5408 5184 5472
rect 5248 5408 5264 5472
rect 5328 5408 5344 5472
rect 5408 5408 5424 5472
rect 5488 5408 5496 5472
rect 5176 5407 5496 5408
rect 9408 5472 9728 5473
rect 9408 5408 9416 5472
rect 9480 5408 9496 5472
rect 9560 5408 9576 5472
rect 9640 5408 9656 5472
rect 9720 5408 9728 5472
rect 9408 5407 9728 5408
rect 3060 4928 3380 4929
rect 3060 4864 3068 4928
rect 3132 4864 3148 4928
rect 3212 4864 3228 4928
rect 3292 4864 3308 4928
rect 3372 4864 3380 4928
rect 3060 4863 3380 4864
rect 7292 4928 7612 4929
rect 7292 4864 7300 4928
rect 7364 4864 7380 4928
rect 7444 4864 7460 4928
rect 7524 4864 7540 4928
rect 7604 4864 7612 4928
rect 7292 4863 7612 4864
rect 11524 4928 11844 4929
rect 11524 4864 11532 4928
rect 11596 4864 11612 4928
rect 11676 4864 11692 4928
rect 11756 4864 11772 4928
rect 11836 4864 11844 4928
rect 11524 4863 11844 4864
rect 5176 4384 5496 4385
rect 5176 4320 5184 4384
rect 5248 4320 5264 4384
rect 5328 4320 5344 4384
rect 5408 4320 5424 4384
rect 5488 4320 5496 4384
rect 5176 4319 5496 4320
rect 9408 4384 9728 4385
rect 9408 4320 9416 4384
rect 9480 4320 9496 4384
rect 9560 4320 9576 4384
rect 9640 4320 9656 4384
rect 9720 4320 9728 4384
rect 9408 4319 9728 4320
rect 3060 3840 3380 3841
rect 3060 3776 3068 3840
rect 3132 3776 3148 3840
rect 3212 3776 3228 3840
rect 3292 3776 3308 3840
rect 3372 3776 3380 3840
rect 3060 3775 3380 3776
rect 7292 3840 7612 3841
rect 7292 3776 7300 3840
rect 7364 3776 7380 3840
rect 7444 3776 7460 3840
rect 7524 3776 7540 3840
rect 7604 3776 7612 3840
rect 7292 3775 7612 3776
rect 11524 3840 11844 3841
rect 11524 3776 11532 3840
rect 11596 3776 11612 3840
rect 11676 3776 11692 3840
rect 11756 3776 11772 3840
rect 11836 3776 11844 3840
rect 11524 3775 11844 3776
rect 13077 3498 13143 3501
rect 14181 3498 14981 3528
rect 13077 3496 14981 3498
rect 13077 3440 13082 3496
rect 13138 3440 14981 3496
rect 13077 3438 14981 3440
rect 13077 3435 13143 3438
rect 14181 3408 14981 3438
rect 5176 3296 5496 3297
rect 5176 3232 5184 3296
rect 5248 3232 5264 3296
rect 5328 3232 5344 3296
rect 5408 3232 5424 3296
rect 5488 3232 5496 3296
rect 5176 3231 5496 3232
rect 9408 3296 9728 3297
rect 9408 3232 9416 3296
rect 9480 3232 9496 3296
rect 9560 3232 9576 3296
rect 9640 3232 9656 3296
rect 9720 3232 9728 3296
rect 9408 3231 9728 3232
rect 0 2818 800 2848
rect 1485 2818 1551 2821
rect 0 2816 1551 2818
rect 0 2760 1490 2816
rect 1546 2760 1551 2816
rect 0 2758 1551 2760
rect 0 2728 800 2758
rect 1485 2755 1551 2758
rect 3060 2752 3380 2753
rect 3060 2688 3068 2752
rect 3132 2688 3148 2752
rect 3212 2688 3228 2752
rect 3292 2688 3308 2752
rect 3372 2688 3380 2752
rect 3060 2687 3380 2688
rect 7292 2752 7612 2753
rect 7292 2688 7300 2752
rect 7364 2688 7380 2752
rect 7444 2688 7460 2752
rect 7524 2688 7540 2752
rect 7604 2688 7612 2752
rect 7292 2687 7612 2688
rect 11524 2752 11844 2753
rect 11524 2688 11532 2752
rect 11596 2688 11612 2752
rect 11676 2688 11692 2752
rect 11756 2688 11772 2752
rect 11836 2688 11844 2752
rect 11524 2687 11844 2688
rect 5176 2208 5496 2209
rect 5176 2144 5184 2208
rect 5248 2144 5264 2208
rect 5328 2144 5344 2208
rect 5408 2144 5424 2208
rect 5488 2144 5496 2208
rect 5176 2143 5496 2144
rect 9408 2208 9728 2209
rect 9408 2144 9416 2208
rect 9480 2144 9496 2208
rect 9560 2144 9576 2208
rect 9640 2144 9656 2208
rect 9720 2144 9728 2208
rect 9408 2143 9728 2144
rect 11973 98 12039 101
rect 14181 98 14981 128
rect 11973 96 14981 98
rect 11973 40 11978 96
rect 12034 40 14981 96
rect 11973 38 14981 40
rect 11973 35 12039 38
rect 14181 8 14981 38
<< via3 >>
rect 3068 14716 3132 14720
rect 3068 14660 3072 14716
rect 3072 14660 3128 14716
rect 3128 14660 3132 14716
rect 3068 14656 3132 14660
rect 3148 14716 3212 14720
rect 3148 14660 3152 14716
rect 3152 14660 3208 14716
rect 3208 14660 3212 14716
rect 3148 14656 3212 14660
rect 3228 14716 3292 14720
rect 3228 14660 3232 14716
rect 3232 14660 3288 14716
rect 3288 14660 3292 14716
rect 3228 14656 3292 14660
rect 3308 14716 3372 14720
rect 3308 14660 3312 14716
rect 3312 14660 3368 14716
rect 3368 14660 3372 14716
rect 3308 14656 3372 14660
rect 7300 14716 7364 14720
rect 7300 14660 7304 14716
rect 7304 14660 7360 14716
rect 7360 14660 7364 14716
rect 7300 14656 7364 14660
rect 7380 14716 7444 14720
rect 7380 14660 7384 14716
rect 7384 14660 7440 14716
rect 7440 14660 7444 14716
rect 7380 14656 7444 14660
rect 7460 14716 7524 14720
rect 7460 14660 7464 14716
rect 7464 14660 7520 14716
rect 7520 14660 7524 14716
rect 7460 14656 7524 14660
rect 7540 14716 7604 14720
rect 7540 14660 7544 14716
rect 7544 14660 7600 14716
rect 7600 14660 7604 14716
rect 7540 14656 7604 14660
rect 11532 14716 11596 14720
rect 11532 14660 11536 14716
rect 11536 14660 11592 14716
rect 11592 14660 11596 14716
rect 11532 14656 11596 14660
rect 11612 14716 11676 14720
rect 11612 14660 11616 14716
rect 11616 14660 11672 14716
rect 11672 14660 11676 14716
rect 11612 14656 11676 14660
rect 11692 14716 11756 14720
rect 11692 14660 11696 14716
rect 11696 14660 11752 14716
rect 11752 14660 11756 14716
rect 11692 14656 11756 14660
rect 11772 14716 11836 14720
rect 11772 14660 11776 14716
rect 11776 14660 11832 14716
rect 11832 14660 11836 14716
rect 11772 14656 11836 14660
rect 5184 14172 5248 14176
rect 5184 14116 5188 14172
rect 5188 14116 5244 14172
rect 5244 14116 5248 14172
rect 5184 14112 5248 14116
rect 5264 14172 5328 14176
rect 5264 14116 5268 14172
rect 5268 14116 5324 14172
rect 5324 14116 5328 14172
rect 5264 14112 5328 14116
rect 5344 14172 5408 14176
rect 5344 14116 5348 14172
rect 5348 14116 5404 14172
rect 5404 14116 5408 14172
rect 5344 14112 5408 14116
rect 5424 14172 5488 14176
rect 5424 14116 5428 14172
rect 5428 14116 5484 14172
rect 5484 14116 5488 14172
rect 5424 14112 5488 14116
rect 9416 14172 9480 14176
rect 9416 14116 9420 14172
rect 9420 14116 9476 14172
rect 9476 14116 9480 14172
rect 9416 14112 9480 14116
rect 9496 14172 9560 14176
rect 9496 14116 9500 14172
rect 9500 14116 9556 14172
rect 9556 14116 9560 14172
rect 9496 14112 9560 14116
rect 9576 14172 9640 14176
rect 9576 14116 9580 14172
rect 9580 14116 9636 14172
rect 9636 14116 9640 14172
rect 9576 14112 9640 14116
rect 9656 14172 9720 14176
rect 9656 14116 9660 14172
rect 9660 14116 9716 14172
rect 9716 14116 9720 14172
rect 9656 14112 9720 14116
rect 3068 13628 3132 13632
rect 3068 13572 3072 13628
rect 3072 13572 3128 13628
rect 3128 13572 3132 13628
rect 3068 13568 3132 13572
rect 3148 13628 3212 13632
rect 3148 13572 3152 13628
rect 3152 13572 3208 13628
rect 3208 13572 3212 13628
rect 3148 13568 3212 13572
rect 3228 13628 3292 13632
rect 3228 13572 3232 13628
rect 3232 13572 3288 13628
rect 3288 13572 3292 13628
rect 3228 13568 3292 13572
rect 3308 13628 3372 13632
rect 3308 13572 3312 13628
rect 3312 13572 3368 13628
rect 3368 13572 3372 13628
rect 3308 13568 3372 13572
rect 7300 13628 7364 13632
rect 7300 13572 7304 13628
rect 7304 13572 7360 13628
rect 7360 13572 7364 13628
rect 7300 13568 7364 13572
rect 7380 13628 7444 13632
rect 7380 13572 7384 13628
rect 7384 13572 7440 13628
rect 7440 13572 7444 13628
rect 7380 13568 7444 13572
rect 7460 13628 7524 13632
rect 7460 13572 7464 13628
rect 7464 13572 7520 13628
rect 7520 13572 7524 13628
rect 7460 13568 7524 13572
rect 7540 13628 7604 13632
rect 7540 13572 7544 13628
rect 7544 13572 7600 13628
rect 7600 13572 7604 13628
rect 7540 13568 7604 13572
rect 11532 13628 11596 13632
rect 11532 13572 11536 13628
rect 11536 13572 11592 13628
rect 11592 13572 11596 13628
rect 11532 13568 11596 13572
rect 11612 13628 11676 13632
rect 11612 13572 11616 13628
rect 11616 13572 11672 13628
rect 11672 13572 11676 13628
rect 11612 13568 11676 13572
rect 11692 13628 11756 13632
rect 11692 13572 11696 13628
rect 11696 13572 11752 13628
rect 11752 13572 11756 13628
rect 11692 13568 11756 13572
rect 11772 13628 11836 13632
rect 11772 13572 11776 13628
rect 11776 13572 11832 13628
rect 11832 13572 11836 13628
rect 11772 13568 11836 13572
rect 5184 13084 5248 13088
rect 5184 13028 5188 13084
rect 5188 13028 5244 13084
rect 5244 13028 5248 13084
rect 5184 13024 5248 13028
rect 5264 13084 5328 13088
rect 5264 13028 5268 13084
rect 5268 13028 5324 13084
rect 5324 13028 5328 13084
rect 5264 13024 5328 13028
rect 5344 13084 5408 13088
rect 5344 13028 5348 13084
rect 5348 13028 5404 13084
rect 5404 13028 5408 13084
rect 5344 13024 5408 13028
rect 5424 13084 5488 13088
rect 5424 13028 5428 13084
rect 5428 13028 5484 13084
rect 5484 13028 5488 13084
rect 5424 13024 5488 13028
rect 9416 13084 9480 13088
rect 9416 13028 9420 13084
rect 9420 13028 9476 13084
rect 9476 13028 9480 13084
rect 9416 13024 9480 13028
rect 9496 13084 9560 13088
rect 9496 13028 9500 13084
rect 9500 13028 9556 13084
rect 9556 13028 9560 13084
rect 9496 13024 9560 13028
rect 9576 13084 9640 13088
rect 9576 13028 9580 13084
rect 9580 13028 9636 13084
rect 9636 13028 9640 13084
rect 9576 13024 9640 13028
rect 9656 13084 9720 13088
rect 9656 13028 9660 13084
rect 9660 13028 9716 13084
rect 9716 13028 9720 13084
rect 9656 13024 9720 13028
rect 3068 12540 3132 12544
rect 3068 12484 3072 12540
rect 3072 12484 3128 12540
rect 3128 12484 3132 12540
rect 3068 12480 3132 12484
rect 3148 12540 3212 12544
rect 3148 12484 3152 12540
rect 3152 12484 3208 12540
rect 3208 12484 3212 12540
rect 3148 12480 3212 12484
rect 3228 12540 3292 12544
rect 3228 12484 3232 12540
rect 3232 12484 3288 12540
rect 3288 12484 3292 12540
rect 3228 12480 3292 12484
rect 3308 12540 3372 12544
rect 3308 12484 3312 12540
rect 3312 12484 3368 12540
rect 3368 12484 3372 12540
rect 3308 12480 3372 12484
rect 7300 12540 7364 12544
rect 7300 12484 7304 12540
rect 7304 12484 7360 12540
rect 7360 12484 7364 12540
rect 7300 12480 7364 12484
rect 7380 12540 7444 12544
rect 7380 12484 7384 12540
rect 7384 12484 7440 12540
rect 7440 12484 7444 12540
rect 7380 12480 7444 12484
rect 7460 12540 7524 12544
rect 7460 12484 7464 12540
rect 7464 12484 7520 12540
rect 7520 12484 7524 12540
rect 7460 12480 7524 12484
rect 7540 12540 7604 12544
rect 7540 12484 7544 12540
rect 7544 12484 7600 12540
rect 7600 12484 7604 12540
rect 7540 12480 7604 12484
rect 11532 12540 11596 12544
rect 11532 12484 11536 12540
rect 11536 12484 11592 12540
rect 11592 12484 11596 12540
rect 11532 12480 11596 12484
rect 11612 12540 11676 12544
rect 11612 12484 11616 12540
rect 11616 12484 11672 12540
rect 11672 12484 11676 12540
rect 11612 12480 11676 12484
rect 11692 12540 11756 12544
rect 11692 12484 11696 12540
rect 11696 12484 11752 12540
rect 11752 12484 11756 12540
rect 11692 12480 11756 12484
rect 11772 12540 11836 12544
rect 11772 12484 11776 12540
rect 11776 12484 11832 12540
rect 11832 12484 11836 12540
rect 11772 12480 11836 12484
rect 5184 11996 5248 12000
rect 5184 11940 5188 11996
rect 5188 11940 5244 11996
rect 5244 11940 5248 11996
rect 5184 11936 5248 11940
rect 5264 11996 5328 12000
rect 5264 11940 5268 11996
rect 5268 11940 5324 11996
rect 5324 11940 5328 11996
rect 5264 11936 5328 11940
rect 5344 11996 5408 12000
rect 5344 11940 5348 11996
rect 5348 11940 5404 11996
rect 5404 11940 5408 11996
rect 5344 11936 5408 11940
rect 5424 11996 5488 12000
rect 5424 11940 5428 11996
rect 5428 11940 5484 11996
rect 5484 11940 5488 11996
rect 5424 11936 5488 11940
rect 9416 11996 9480 12000
rect 9416 11940 9420 11996
rect 9420 11940 9476 11996
rect 9476 11940 9480 11996
rect 9416 11936 9480 11940
rect 9496 11996 9560 12000
rect 9496 11940 9500 11996
rect 9500 11940 9556 11996
rect 9556 11940 9560 11996
rect 9496 11936 9560 11940
rect 9576 11996 9640 12000
rect 9576 11940 9580 11996
rect 9580 11940 9636 11996
rect 9636 11940 9640 11996
rect 9576 11936 9640 11940
rect 9656 11996 9720 12000
rect 9656 11940 9660 11996
rect 9660 11940 9716 11996
rect 9716 11940 9720 11996
rect 9656 11936 9720 11940
rect 3068 11452 3132 11456
rect 3068 11396 3072 11452
rect 3072 11396 3128 11452
rect 3128 11396 3132 11452
rect 3068 11392 3132 11396
rect 3148 11452 3212 11456
rect 3148 11396 3152 11452
rect 3152 11396 3208 11452
rect 3208 11396 3212 11452
rect 3148 11392 3212 11396
rect 3228 11452 3292 11456
rect 3228 11396 3232 11452
rect 3232 11396 3288 11452
rect 3288 11396 3292 11452
rect 3228 11392 3292 11396
rect 3308 11452 3372 11456
rect 3308 11396 3312 11452
rect 3312 11396 3368 11452
rect 3368 11396 3372 11452
rect 3308 11392 3372 11396
rect 7300 11452 7364 11456
rect 7300 11396 7304 11452
rect 7304 11396 7360 11452
rect 7360 11396 7364 11452
rect 7300 11392 7364 11396
rect 7380 11452 7444 11456
rect 7380 11396 7384 11452
rect 7384 11396 7440 11452
rect 7440 11396 7444 11452
rect 7380 11392 7444 11396
rect 7460 11452 7524 11456
rect 7460 11396 7464 11452
rect 7464 11396 7520 11452
rect 7520 11396 7524 11452
rect 7460 11392 7524 11396
rect 7540 11452 7604 11456
rect 7540 11396 7544 11452
rect 7544 11396 7600 11452
rect 7600 11396 7604 11452
rect 7540 11392 7604 11396
rect 11532 11452 11596 11456
rect 11532 11396 11536 11452
rect 11536 11396 11592 11452
rect 11592 11396 11596 11452
rect 11532 11392 11596 11396
rect 11612 11452 11676 11456
rect 11612 11396 11616 11452
rect 11616 11396 11672 11452
rect 11672 11396 11676 11452
rect 11612 11392 11676 11396
rect 11692 11452 11756 11456
rect 11692 11396 11696 11452
rect 11696 11396 11752 11452
rect 11752 11396 11756 11452
rect 11692 11392 11756 11396
rect 11772 11452 11836 11456
rect 11772 11396 11776 11452
rect 11776 11396 11832 11452
rect 11832 11396 11836 11452
rect 11772 11392 11836 11396
rect 5184 10908 5248 10912
rect 5184 10852 5188 10908
rect 5188 10852 5244 10908
rect 5244 10852 5248 10908
rect 5184 10848 5248 10852
rect 5264 10908 5328 10912
rect 5264 10852 5268 10908
rect 5268 10852 5324 10908
rect 5324 10852 5328 10908
rect 5264 10848 5328 10852
rect 5344 10908 5408 10912
rect 5344 10852 5348 10908
rect 5348 10852 5404 10908
rect 5404 10852 5408 10908
rect 5344 10848 5408 10852
rect 5424 10908 5488 10912
rect 5424 10852 5428 10908
rect 5428 10852 5484 10908
rect 5484 10852 5488 10908
rect 5424 10848 5488 10852
rect 9416 10908 9480 10912
rect 9416 10852 9420 10908
rect 9420 10852 9476 10908
rect 9476 10852 9480 10908
rect 9416 10848 9480 10852
rect 9496 10908 9560 10912
rect 9496 10852 9500 10908
rect 9500 10852 9556 10908
rect 9556 10852 9560 10908
rect 9496 10848 9560 10852
rect 9576 10908 9640 10912
rect 9576 10852 9580 10908
rect 9580 10852 9636 10908
rect 9636 10852 9640 10908
rect 9576 10848 9640 10852
rect 9656 10908 9720 10912
rect 9656 10852 9660 10908
rect 9660 10852 9716 10908
rect 9716 10852 9720 10908
rect 9656 10848 9720 10852
rect 3068 10364 3132 10368
rect 3068 10308 3072 10364
rect 3072 10308 3128 10364
rect 3128 10308 3132 10364
rect 3068 10304 3132 10308
rect 3148 10364 3212 10368
rect 3148 10308 3152 10364
rect 3152 10308 3208 10364
rect 3208 10308 3212 10364
rect 3148 10304 3212 10308
rect 3228 10364 3292 10368
rect 3228 10308 3232 10364
rect 3232 10308 3288 10364
rect 3288 10308 3292 10364
rect 3228 10304 3292 10308
rect 3308 10364 3372 10368
rect 3308 10308 3312 10364
rect 3312 10308 3368 10364
rect 3368 10308 3372 10364
rect 3308 10304 3372 10308
rect 7300 10364 7364 10368
rect 7300 10308 7304 10364
rect 7304 10308 7360 10364
rect 7360 10308 7364 10364
rect 7300 10304 7364 10308
rect 7380 10364 7444 10368
rect 7380 10308 7384 10364
rect 7384 10308 7440 10364
rect 7440 10308 7444 10364
rect 7380 10304 7444 10308
rect 7460 10364 7524 10368
rect 7460 10308 7464 10364
rect 7464 10308 7520 10364
rect 7520 10308 7524 10364
rect 7460 10304 7524 10308
rect 7540 10364 7604 10368
rect 7540 10308 7544 10364
rect 7544 10308 7600 10364
rect 7600 10308 7604 10364
rect 7540 10304 7604 10308
rect 11532 10364 11596 10368
rect 11532 10308 11536 10364
rect 11536 10308 11592 10364
rect 11592 10308 11596 10364
rect 11532 10304 11596 10308
rect 11612 10364 11676 10368
rect 11612 10308 11616 10364
rect 11616 10308 11672 10364
rect 11672 10308 11676 10364
rect 11612 10304 11676 10308
rect 11692 10364 11756 10368
rect 11692 10308 11696 10364
rect 11696 10308 11752 10364
rect 11752 10308 11756 10364
rect 11692 10304 11756 10308
rect 11772 10364 11836 10368
rect 11772 10308 11776 10364
rect 11776 10308 11832 10364
rect 11832 10308 11836 10364
rect 11772 10304 11836 10308
rect 5184 9820 5248 9824
rect 5184 9764 5188 9820
rect 5188 9764 5244 9820
rect 5244 9764 5248 9820
rect 5184 9760 5248 9764
rect 5264 9820 5328 9824
rect 5264 9764 5268 9820
rect 5268 9764 5324 9820
rect 5324 9764 5328 9820
rect 5264 9760 5328 9764
rect 5344 9820 5408 9824
rect 5344 9764 5348 9820
rect 5348 9764 5404 9820
rect 5404 9764 5408 9820
rect 5344 9760 5408 9764
rect 5424 9820 5488 9824
rect 5424 9764 5428 9820
rect 5428 9764 5484 9820
rect 5484 9764 5488 9820
rect 5424 9760 5488 9764
rect 9416 9820 9480 9824
rect 9416 9764 9420 9820
rect 9420 9764 9476 9820
rect 9476 9764 9480 9820
rect 9416 9760 9480 9764
rect 9496 9820 9560 9824
rect 9496 9764 9500 9820
rect 9500 9764 9556 9820
rect 9556 9764 9560 9820
rect 9496 9760 9560 9764
rect 9576 9820 9640 9824
rect 9576 9764 9580 9820
rect 9580 9764 9636 9820
rect 9636 9764 9640 9820
rect 9576 9760 9640 9764
rect 9656 9820 9720 9824
rect 9656 9764 9660 9820
rect 9660 9764 9716 9820
rect 9716 9764 9720 9820
rect 9656 9760 9720 9764
rect 3068 9276 3132 9280
rect 3068 9220 3072 9276
rect 3072 9220 3128 9276
rect 3128 9220 3132 9276
rect 3068 9216 3132 9220
rect 3148 9276 3212 9280
rect 3148 9220 3152 9276
rect 3152 9220 3208 9276
rect 3208 9220 3212 9276
rect 3148 9216 3212 9220
rect 3228 9276 3292 9280
rect 3228 9220 3232 9276
rect 3232 9220 3288 9276
rect 3288 9220 3292 9276
rect 3228 9216 3292 9220
rect 3308 9276 3372 9280
rect 3308 9220 3312 9276
rect 3312 9220 3368 9276
rect 3368 9220 3372 9276
rect 3308 9216 3372 9220
rect 7300 9276 7364 9280
rect 7300 9220 7304 9276
rect 7304 9220 7360 9276
rect 7360 9220 7364 9276
rect 7300 9216 7364 9220
rect 7380 9276 7444 9280
rect 7380 9220 7384 9276
rect 7384 9220 7440 9276
rect 7440 9220 7444 9276
rect 7380 9216 7444 9220
rect 7460 9276 7524 9280
rect 7460 9220 7464 9276
rect 7464 9220 7520 9276
rect 7520 9220 7524 9276
rect 7460 9216 7524 9220
rect 7540 9276 7604 9280
rect 7540 9220 7544 9276
rect 7544 9220 7600 9276
rect 7600 9220 7604 9276
rect 7540 9216 7604 9220
rect 11532 9276 11596 9280
rect 11532 9220 11536 9276
rect 11536 9220 11592 9276
rect 11592 9220 11596 9276
rect 11532 9216 11596 9220
rect 11612 9276 11676 9280
rect 11612 9220 11616 9276
rect 11616 9220 11672 9276
rect 11672 9220 11676 9276
rect 11612 9216 11676 9220
rect 11692 9276 11756 9280
rect 11692 9220 11696 9276
rect 11696 9220 11752 9276
rect 11752 9220 11756 9276
rect 11692 9216 11756 9220
rect 11772 9276 11836 9280
rect 11772 9220 11776 9276
rect 11776 9220 11832 9276
rect 11832 9220 11836 9276
rect 11772 9216 11836 9220
rect 5184 8732 5248 8736
rect 5184 8676 5188 8732
rect 5188 8676 5244 8732
rect 5244 8676 5248 8732
rect 5184 8672 5248 8676
rect 5264 8732 5328 8736
rect 5264 8676 5268 8732
rect 5268 8676 5324 8732
rect 5324 8676 5328 8732
rect 5264 8672 5328 8676
rect 5344 8732 5408 8736
rect 5344 8676 5348 8732
rect 5348 8676 5404 8732
rect 5404 8676 5408 8732
rect 5344 8672 5408 8676
rect 5424 8732 5488 8736
rect 5424 8676 5428 8732
rect 5428 8676 5484 8732
rect 5484 8676 5488 8732
rect 5424 8672 5488 8676
rect 9416 8732 9480 8736
rect 9416 8676 9420 8732
rect 9420 8676 9476 8732
rect 9476 8676 9480 8732
rect 9416 8672 9480 8676
rect 9496 8732 9560 8736
rect 9496 8676 9500 8732
rect 9500 8676 9556 8732
rect 9556 8676 9560 8732
rect 9496 8672 9560 8676
rect 9576 8732 9640 8736
rect 9576 8676 9580 8732
rect 9580 8676 9636 8732
rect 9636 8676 9640 8732
rect 9576 8672 9640 8676
rect 9656 8732 9720 8736
rect 9656 8676 9660 8732
rect 9660 8676 9716 8732
rect 9716 8676 9720 8732
rect 9656 8672 9720 8676
rect 3068 8188 3132 8192
rect 3068 8132 3072 8188
rect 3072 8132 3128 8188
rect 3128 8132 3132 8188
rect 3068 8128 3132 8132
rect 3148 8188 3212 8192
rect 3148 8132 3152 8188
rect 3152 8132 3208 8188
rect 3208 8132 3212 8188
rect 3148 8128 3212 8132
rect 3228 8188 3292 8192
rect 3228 8132 3232 8188
rect 3232 8132 3288 8188
rect 3288 8132 3292 8188
rect 3228 8128 3292 8132
rect 3308 8188 3372 8192
rect 3308 8132 3312 8188
rect 3312 8132 3368 8188
rect 3368 8132 3372 8188
rect 3308 8128 3372 8132
rect 7300 8188 7364 8192
rect 7300 8132 7304 8188
rect 7304 8132 7360 8188
rect 7360 8132 7364 8188
rect 7300 8128 7364 8132
rect 7380 8188 7444 8192
rect 7380 8132 7384 8188
rect 7384 8132 7440 8188
rect 7440 8132 7444 8188
rect 7380 8128 7444 8132
rect 7460 8188 7524 8192
rect 7460 8132 7464 8188
rect 7464 8132 7520 8188
rect 7520 8132 7524 8188
rect 7460 8128 7524 8132
rect 7540 8188 7604 8192
rect 7540 8132 7544 8188
rect 7544 8132 7600 8188
rect 7600 8132 7604 8188
rect 7540 8128 7604 8132
rect 11532 8188 11596 8192
rect 11532 8132 11536 8188
rect 11536 8132 11592 8188
rect 11592 8132 11596 8188
rect 11532 8128 11596 8132
rect 11612 8188 11676 8192
rect 11612 8132 11616 8188
rect 11616 8132 11672 8188
rect 11672 8132 11676 8188
rect 11612 8128 11676 8132
rect 11692 8188 11756 8192
rect 11692 8132 11696 8188
rect 11696 8132 11752 8188
rect 11752 8132 11756 8188
rect 11692 8128 11756 8132
rect 11772 8188 11836 8192
rect 11772 8132 11776 8188
rect 11776 8132 11832 8188
rect 11832 8132 11836 8188
rect 11772 8128 11836 8132
rect 5184 7644 5248 7648
rect 5184 7588 5188 7644
rect 5188 7588 5244 7644
rect 5244 7588 5248 7644
rect 5184 7584 5248 7588
rect 5264 7644 5328 7648
rect 5264 7588 5268 7644
rect 5268 7588 5324 7644
rect 5324 7588 5328 7644
rect 5264 7584 5328 7588
rect 5344 7644 5408 7648
rect 5344 7588 5348 7644
rect 5348 7588 5404 7644
rect 5404 7588 5408 7644
rect 5344 7584 5408 7588
rect 5424 7644 5488 7648
rect 5424 7588 5428 7644
rect 5428 7588 5484 7644
rect 5484 7588 5488 7644
rect 5424 7584 5488 7588
rect 9416 7644 9480 7648
rect 9416 7588 9420 7644
rect 9420 7588 9476 7644
rect 9476 7588 9480 7644
rect 9416 7584 9480 7588
rect 9496 7644 9560 7648
rect 9496 7588 9500 7644
rect 9500 7588 9556 7644
rect 9556 7588 9560 7644
rect 9496 7584 9560 7588
rect 9576 7644 9640 7648
rect 9576 7588 9580 7644
rect 9580 7588 9636 7644
rect 9636 7588 9640 7644
rect 9576 7584 9640 7588
rect 9656 7644 9720 7648
rect 9656 7588 9660 7644
rect 9660 7588 9716 7644
rect 9716 7588 9720 7644
rect 9656 7584 9720 7588
rect 3068 7100 3132 7104
rect 3068 7044 3072 7100
rect 3072 7044 3128 7100
rect 3128 7044 3132 7100
rect 3068 7040 3132 7044
rect 3148 7100 3212 7104
rect 3148 7044 3152 7100
rect 3152 7044 3208 7100
rect 3208 7044 3212 7100
rect 3148 7040 3212 7044
rect 3228 7100 3292 7104
rect 3228 7044 3232 7100
rect 3232 7044 3288 7100
rect 3288 7044 3292 7100
rect 3228 7040 3292 7044
rect 3308 7100 3372 7104
rect 3308 7044 3312 7100
rect 3312 7044 3368 7100
rect 3368 7044 3372 7100
rect 3308 7040 3372 7044
rect 7300 7100 7364 7104
rect 7300 7044 7304 7100
rect 7304 7044 7360 7100
rect 7360 7044 7364 7100
rect 7300 7040 7364 7044
rect 7380 7100 7444 7104
rect 7380 7044 7384 7100
rect 7384 7044 7440 7100
rect 7440 7044 7444 7100
rect 7380 7040 7444 7044
rect 7460 7100 7524 7104
rect 7460 7044 7464 7100
rect 7464 7044 7520 7100
rect 7520 7044 7524 7100
rect 7460 7040 7524 7044
rect 7540 7100 7604 7104
rect 7540 7044 7544 7100
rect 7544 7044 7600 7100
rect 7600 7044 7604 7100
rect 7540 7040 7604 7044
rect 11532 7100 11596 7104
rect 11532 7044 11536 7100
rect 11536 7044 11592 7100
rect 11592 7044 11596 7100
rect 11532 7040 11596 7044
rect 11612 7100 11676 7104
rect 11612 7044 11616 7100
rect 11616 7044 11672 7100
rect 11672 7044 11676 7100
rect 11612 7040 11676 7044
rect 11692 7100 11756 7104
rect 11692 7044 11696 7100
rect 11696 7044 11752 7100
rect 11752 7044 11756 7100
rect 11692 7040 11756 7044
rect 11772 7100 11836 7104
rect 11772 7044 11776 7100
rect 11776 7044 11832 7100
rect 11832 7044 11836 7100
rect 11772 7040 11836 7044
rect 5184 6556 5248 6560
rect 5184 6500 5188 6556
rect 5188 6500 5244 6556
rect 5244 6500 5248 6556
rect 5184 6496 5248 6500
rect 5264 6556 5328 6560
rect 5264 6500 5268 6556
rect 5268 6500 5324 6556
rect 5324 6500 5328 6556
rect 5264 6496 5328 6500
rect 5344 6556 5408 6560
rect 5344 6500 5348 6556
rect 5348 6500 5404 6556
rect 5404 6500 5408 6556
rect 5344 6496 5408 6500
rect 5424 6556 5488 6560
rect 5424 6500 5428 6556
rect 5428 6500 5484 6556
rect 5484 6500 5488 6556
rect 5424 6496 5488 6500
rect 9416 6556 9480 6560
rect 9416 6500 9420 6556
rect 9420 6500 9476 6556
rect 9476 6500 9480 6556
rect 9416 6496 9480 6500
rect 9496 6556 9560 6560
rect 9496 6500 9500 6556
rect 9500 6500 9556 6556
rect 9556 6500 9560 6556
rect 9496 6496 9560 6500
rect 9576 6556 9640 6560
rect 9576 6500 9580 6556
rect 9580 6500 9636 6556
rect 9636 6500 9640 6556
rect 9576 6496 9640 6500
rect 9656 6556 9720 6560
rect 9656 6500 9660 6556
rect 9660 6500 9716 6556
rect 9716 6500 9720 6556
rect 9656 6496 9720 6500
rect 3068 6012 3132 6016
rect 3068 5956 3072 6012
rect 3072 5956 3128 6012
rect 3128 5956 3132 6012
rect 3068 5952 3132 5956
rect 3148 6012 3212 6016
rect 3148 5956 3152 6012
rect 3152 5956 3208 6012
rect 3208 5956 3212 6012
rect 3148 5952 3212 5956
rect 3228 6012 3292 6016
rect 3228 5956 3232 6012
rect 3232 5956 3288 6012
rect 3288 5956 3292 6012
rect 3228 5952 3292 5956
rect 3308 6012 3372 6016
rect 3308 5956 3312 6012
rect 3312 5956 3368 6012
rect 3368 5956 3372 6012
rect 3308 5952 3372 5956
rect 7300 6012 7364 6016
rect 7300 5956 7304 6012
rect 7304 5956 7360 6012
rect 7360 5956 7364 6012
rect 7300 5952 7364 5956
rect 7380 6012 7444 6016
rect 7380 5956 7384 6012
rect 7384 5956 7440 6012
rect 7440 5956 7444 6012
rect 7380 5952 7444 5956
rect 7460 6012 7524 6016
rect 7460 5956 7464 6012
rect 7464 5956 7520 6012
rect 7520 5956 7524 6012
rect 7460 5952 7524 5956
rect 7540 6012 7604 6016
rect 7540 5956 7544 6012
rect 7544 5956 7600 6012
rect 7600 5956 7604 6012
rect 7540 5952 7604 5956
rect 11532 6012 11596 6016
rect 11532 5956 11536 6012
rect 11536 5956 11592 6012
rect 11592 5956 11596 6012
rect 11532 5952 11596 5956
rect 11612 6012 11676 6016
rect 11612 5956 11616 6012
rect 11616 5956 11672 6012
rect 11672 5956 11676 6012
rect 11612 5952 11676 5956
rect 11692 6012 11756 6016
rect 11692 5956 11696 6012
rect 11696 5956 11752 6012
rect 11752 5956 11756 6012
rect 11692 5952 11756 5956
rect 11772 6012 11836 6016
rect 11772 5956 11776 6012
rect 11776 5956 11832 6012
rect 11832 5956 11836 6012
rect 11772 5952 11836 5956
rect 5184 5468 5248 5472
rect 5184 5412 5188 5468
rect 5188 5412 5244 5468
rect 5244 5412 5248 5468
rect 5184 5408 5248 5412
rect 5264 5468 5328 5472
rect 5264 5412 5268 5468
rect 5268 5412 5324 5468
rect 5324 5412 5328 5468
rect 5264 5408 5328 5412
rect 5344 5468 5408 5472
rect 5344 5412 5348 5468
rect 5348 5412 5404 5468
rect 5404 5412 5408 5468
rect 5344 5408 5408 5412
rect 5424 5468 5488 5472
rect 5424 5412 5428 5468
rect 5428 5412 5484 5468
rect 5484 5412 5488 5468
rect 5424 5408 5488 5412
rect 9416 5468 9480 5472
rect 9416 5412 9420 5468
rect 9420 5412 9476 5468
rect 9476 5412 9480 5468
rect 9416 5408 9480 5412
rect 9496 5468 9560 5472
rect 9496 5412 9500 5468
rect 9500 5412 9556 5468
rect 9556 5412 9560 5468
rect 9496 5408 9560 5412
rect 9576 5468 9640 5472
rect 9576 5412 9580 5468
rect 9580 5412 9636 5468
rect 9636 5412 9640 5468
rect 9576 5408 9640 5412
rect 9656 5468 9720 5472
rect 9656 5412 9660 5468
rect 9660 5412 9716 5468
rect 9716 5412 9720 5468
rect 9656 5408 9720 5412
rect 3068 4924 3132 4928
rect 3068 4868 3072 4924
rect 3072 4868 3128 4924
rect 3128 4868 3132 4924
rect 3068 4864 3132 4868
rect 3148 4924 3212 4928
rect 3148 4868 3152 4924
rect 3152 4868 3208 4924
rect 3208 4868 3212 4924
rect 3148 4864 3212 4868
rect 3228 4924 3292 4928
rect 3228 4868 3232 4924
rect 3232 4868 3288 4924
rect 3288 4868 3292 4924
rect 3228 4864 3292 4868
rect 3308 4924 3372 4928
rect 3308 4868 3312 4924
rect 3312 4868 3368 4924
rect 3368 4868 3372 4924
rect 3308 4864 3372 4868
rect 7300 4924 7364 4928
rect 7300 4868 7304 4924
rect 7304 4868 7360 4924
rect 7360 4868 7364 4924
rect 7300 4864 7364 4868
rect 7380 4924 7444 4928
rect 7380 4868 7384 4924
rect 7384 4868 7440 4924
rect 7440 4868 7444 4924
rect 7380 4864 7444 4868
rect 7460 4924 7524 4928
rect 7460 4868 7464 4924
rect 7464 4868 7520 4924
rect 7520 4868 7524 4924
rect 7460 4864 7524 4868
rect 7540 4924 7604 4928
rect 7540 4868 7544 4924
rect 7544 4868 7600 4924
rect 7600 4868 7604 4924
rect 7540 4864 7604 4868
rect 11532 4924 11596 4928
rect 11532 4868 11536 4924
rect 11536 4868 11592 4924
rect 11592 4868 11596 4924
rect 11532 4864 11596 4868
rect 11612 4924 11676 4928
rect 11612 4868 11616 4924
rect 11616 4868 11672 4924
rect 11672 4868 11676 4924
rect 11612 4864 11676 4868
rect 11692 4924 11756 4928
rect 11692 4868 11696 4924
rect 11696 4868 11752 4924
rect 11752 4868 11756 4924
rect 11692 4864 11756 4868
rect 11772 4924 11836 4928
rect 11772 4868 11776 4924
rect 11776 4868 11832 4924
rect 11832 4868 11836 4924
rect 11772 4864 11836 4868
rect 5184 4380 5248 4384
rect 5184 4324 5188 4380
rect 5188 4324 5244 4380
rect 5244 4324 5248 4380
rect 5184 4320 5248 4324
rect 5264 4380 5328 4384
rect 5264 4324 5268 4380
rect 5268 4324 5324 4380
rect 5324 4324 5328 4380
rect 5264 4320 5328 4324
rect 5344 4380 5408 4384
rect 5344 4324 5348 4380
rect 5348 4324 5404 4380
rect 5404 4324 5408 4380
rect 5344 4320 5408 4324
rect 5424 4380 5488 4384
rect 5424 4324 5428 4380
rect 5428 4324 5484 4380
rect 5484 4324 5488 4380
rect 5424 4320 5488 4324
rect 9416 4380 9480 4384
rect 9416 4324 9420 4380
rect 9420 4324 9476 4380
rect 9476 4324 9480 4380
rect 9416 4320 9480 4324
rect 9496 4380 9560 4384
rect 9496 4324 9500 4380
rect 9500 4324 9556 4380
rect 9556 4324 9560 4380
rect 9496 4320 9560 4324
rect 9576 4380 9640 4384
rect 9576 4324 9580 4380
rect 9580 4324 9636 4380
rect 9636 4324 9640 4380
rect 9576 4320 9640 4324
rect 9656 4380 9720 4384
rect 9656 4324 9660 4380
rect 9660 4324 9716 4380
rect 9716 4324 9720 4380
rect 9656 4320 9720 4324
rect 3068 3836 3132 3840
rect 3068 3780 3072 3836
rect 3072 3780 3128 3836
rect 3128 3780 3132 3836
rect 3068 3776 3132 3780
rect 3148 3836 3212 3840
rect 3148 3780 3152 3836
rect 3152 3780 3208 3836
rect 3208 3780 3212 3836
rect 3148 3776 3212 3780
rect 3228 3836 3292 3840
rect 3228 3780 3232 3836
rect 3232 3780 3288 3836
rect 3288 3780 3292 3836
rect 3228 3776 3292 3780
rect 3308 3836 3372 3840
rect 3308 3780 3312 3836
rect 3312 3780 3368 3836
rect 3368 3780 3372 3836
rect 3308 3776 3372 3780
rect 7300 3836 7364 3840
rect 7300 3780 7304 3836
rect 7304 3780 7360 3836
rect 7360 3780 7364 3836
rect 7300 3776 7364 3780
rect 7380 3836 7444 3840
rect 7380 3780 7384 3836
rect 7384 3780 7440 3836
rect 7440 3780 7444 3836
rect 7380 3776 7444 3780
rect 7460 3836 7524 3840
rect 7460 3780 7464 3836
rect 7464 3780 7520 3836
rect 7520 3780 7524 3836
rect 7460 3776 7524 3780
rect 7540 3836 7604 3840
rect 7540 3780 7544 3836
rect 7544 3780 7600 3836
rect 7600 3780 7604 3836
rect 7540 3776 7604 3780
rect 11532 3836 11596 3840
rect 11532 3780 11536 3836
rect 11536 3780 11592 3836
rect 11592 3780 11596 3836
rect 11532 3776 11596 3780
rect 11612 3836 11676 3840
rect 11612 3780 11616 3836
rect 11616 3780 11672 3836
rect 11672 3780 11676 3836
rect 11612 3776 11676 3780
rect 11692 3836 11756 3840
rect 11692 3780 11696 3836
rect 11696 3780 11752 3836
rect 11752 3780 11756 3836
rect 11692 3776 11756 3780
rect 11772 3836 11836 3840
rect 11772 3780 11776 3836
rect 11776 3780 11832 3836
rect 11832 3780 11836 3836
rect 11772 3776 11836 3780
rect 5184 3292 5248 3296
rect 5184 3236 5188 3292
rect 5188 3236 5244 3292
rect 5244 3236 5248 3292
rect 5184 3232 5248 3236
rect 5264 3292 5328 3296
rect 5264 3236 5268 3292
rect 5268 3236 5324 3292
rect 5324 3236 5328 3292
rect 5264 3232 5328 3236
rect 5344 3292 5408 3296
rect 5344 3236 5348 3292
rect 5348 3236 5404 3292
rect 5404 3236 5408 3292
rect 5344 3232 5408 3236
rect 5424 3292 5488 3296
rect 5424 3236 5428 3292
rect 5428 3236 5484 3292
rect 5484 3236 5488 3292
rect 5424 3232 5488 3236
rect 9416 3292 9480 3296
rect 9416 3236 9420 3292
rect 9420 3236 9476 3292
rect 9476 3236 9480 3292
rect 9416 3232 9480 3236
rect 9496 3292 9560 3296
rect 9496 3236 9500 3292
rect 9500 3236 9556 3292
rect 9556 3236 9560 3292
rect 9496 3232 9560 3236
rect 9576 3292 9640 3296
rect 9576 3236 9580 3292
rect 9580 3236 9636 3292
rect 9636 3236 9640 3292
rect 9576 3232 9640 3236
rect 9656 3292 9720 3296
rect 9656 3236 9660 3292
rect 9660 3236 9716 3292
rect 9716 3236 9720 3292
rect 9656 3232 9720 3236
rect 3068 2748 3132 2752
rect 3068 2692 3072 2748
rect 3072 2692 3128 2748
rect 3128 2692 3132 2748
rect 3068 2688 3132 2692
rect 3148 2748 3212 2752
rect 3148 2692 3152 2748
rect 3152 2692 3208 2748
rect 3208 2692 3212 2748
rect 3148 2688 3212 2692
rect 3228 2748 3292 2752
rect 3228 2692 3232 2748
rect 3232 2692 3288 2748
rect 3288 2692 3292 2748
rect 3228 2688 3292 2692
rect 3308 2748 3372 2752
rect 3308 2692 3312 2748
rect 3312 2692 3368 2748
rect 3368 2692 3372 2748
rect 3308 2688 3372 2692
rect 7300 2748 7364 2752
rect 7300 2692 7304 2748
rect 7304 2692 7360 2748
rect 7360 2692 7364 2748
rect 7300 2688 7364 2692
rect 7380 2748 7444 2752
rect 7380 2692 7384 2748
rect 7384 2692 7440 2748
rect 7440 2692 7444 2748
rect 7380 2688 7444 2692
rect 7460 2748 7524 2752
rect 7460 2692 7464 2748
rect 7464 2692 7520 2748
rect 7520 2692 7524 2748
rect 7460 2688 7524 2692
rect 7540 2748 7604 2752
rect 7540 2692 7544 2748
rect 7544 2692 7600 2748
rect 7600 2692 7604 2748
rect 7540 2688 7604 2692
rect 11532 2748 11596 2752
rect 11532 2692 11536 2748
rect 11536 2692 11592 2748
rect 11592 2692 11596 2748
rect 11532 2688 11596 2692
rect 11612 2748 11676 2752
rect 11612 2692 11616 2748
rect 11616 2692 11672 2748
rect 11672 2692 11676 2748
rect 11612 2688 11676 2692
rect 11692 2748 11756 2752
rect 11692 2692 11696 2748
rect 11696 2692 11752 2748
rect 11752 2692 11756 2748
rect 11692 2688 11756 2692
rect 11772 2748 11836 2752
rect 11772 2692 11776 2748
rect 11776 2692 11832 2748
rect 11832 2692 11836 2748
rect 11772 2688 11836 2692
rect 5184 2204 5248 2208
rect 5184 2148 5188 2204
rect 5188 2148 5244 2204
rect 5244 2148 5248 2204
rect 5184 2144 5248 2148
rect 5264 2204 5328 2208
rect 5264 2148 5268 2204
rect 5268 2148 5324 2204
rect 5324 2148 5328 2204
rect 5264 2144 5328 2148
rect 5344 2204 5408 2208
rect 5344 2148 5348 2204
rect 5348 2148 5404 2204
rect 5404 2148 5408 2204
rect 5344 2144 5408 2148
rect 5424 2204 5488 2208
rect 5424 2148 5428 2204
rect 5428 2148 5484 2204
rect 5484 2148 5488 2204
rect 5424 2144 5488 2148
rect 9416 2204 9480 2208
rect 9416 2148 9420 2204
rect 9420 2148 9476 2204
rect 9476 2148 9480 2204
rect 9416 2144 9480 2148
rect 9496 2204 9560 2208
rect 9496 2148 9500 2204
rect 9500 2148 9556 2204
rect 9556 2148 9560 2204
rect 9496 2144 9560 2148
rect 9576 2204 9640 2208
rect 9576 2148 9580 2204
rect 9580 2148 9636 2204
rect 9636 2148 9640 2204
rect 9576 2144 9640 2148
rect 9656 2204 9720 2208
rect 9656 2148 9660 2204
rect 9660 2148 9716 2204
rect 9716 2148 9720 2204
rect 9656 2144 9720 2148
<< metal4 >>
rect 3060 14720 3380 14736
rect 3060 14656 3068 14720
rect 3132 14656 3148 14720
rect 3212 14656 3228 14720
rect 3292 14656 3308 14720
rect 3372 14656 3380 14720
rect 3060 13632 3380 14656
rect 3060 13568 3068 13632
rect 3132 13568 3148 13632
rect 3212 13568 3228 13632
rect 3292 13568 3308 13632
rect 3372 13568 3380 13632
rect 3060 12672 3380 13568
rect 3060 12544 3102 12672
rect 3338 12544 3380 12672
rect 3060 12480 3068 12544
rect 3372 12480 3380 12544
rect 3060 12436 3102 12480
rect 3338 12436 3380 12480
rect 3060 11456 3380 12436
rect 3060 11392 3068 11456
rect 3132 11392 3148 11456
rect 3212 11392 3228 11456
rect 3292 11392 3308 11456
rect 3372 11392 3380 11456
rect 3060 10368 3380 11392
rect 3060 10304 3068 10368
rect 3132 10304 3148 10368
rect 3212 10304 3228 10368
rect 3292 10304 3308 10368
rect 3372 10304 3380 10368
rect 3060 9280 3380 10304
rect 3060 9216 3068 9280
rect 3132 9216 3148 9280
rect 3212 9216 3228 9280
rect 3292 9216 3308 9280
rect 3372 9216 3380 9280
rect 3060 8502 3380 9216
rect 3060 8266 3102 8502
rect 3338 8266 3380 8502
rect 3060 8192 3380 8266
rect 3060 8128 3068 8192
rect 3132 8128 3148 8192
rect 3212 8128 3228 8192
rect 3292 8128 3308 8192
rect 3372 8128 3380 8192
rect 3060 7104 3380 8128
rect 3060 7040 3068 7104
rect 3132 7040 3148 7104
rect 3212 7040 3228 7104
rect 3292 7040 3308 7104
rect 3372 7040 3380 7104
rect 3060 6016 3380 7040
rect 3060 5952 3068 6016
rect 3132 5952 3148 6016
rect 3212 5952 3228 6016
rect 3292 5952 3308 6016
rect 3372 5952 3380 6016
rect 3060 4928 3380 5952
rect 3060 4864 3068 4928
rect 3132 4864 3148 4928
rect 3212 4864 3228 4928
rect 3292 4864 3308 4928
rect 3372 4864 3380 4928
rect 3060 4331 3380 4864
rect 3060 4095 3102 4331
rect 3338 4095 3380 4331
rect 3060 3840 3380 4095
rect 3060 3776 3068 3840
rect 3132 3776 3148 3840
rect 3212 3776 3228 3840
rect 3292 3776 3308 3840
rect 3372 3776 3380 3840
rect 3060 2752 3380 3776
rect 3060 2688 3068 2752
rect 3132 2688 3148 2752
rect 3212 2688 3228 2752
rect 3292 2688 3308 2752
rect 3372 2688 3380 2752
rect 3060 2128 3380 2688
rect 5176 14176 5496 14736
rect 5176 14112 5184 14176
rect 5248 14112 5264 14176
rect 5328 14112 5344 14176
rect 5408 14112 5424 14176
rect 5488 14112 5496 14176
rect 5176 13088 5496 14112
rect 5176 13024 5184 13088
rect 5248 13024 5264 13088
rect 5328 13024 5344 13088
rect 5408 13024 5424 13088
rect 5488 13024 5496 13088
rect 5176 12000 5496 13024
rect 5176 11936 5184 12000
rect 5248 11936 5264 12000
rect 5328 11936 5344 12000
rect 5408 11936 5424 12000
rect 5488 11936 5496 12000
rect 5176 10912 5496 11936
rect 5176 10848 5184 10912
rect 5248 10848 5264 10912
rect 5328 10848 5344 10912
rect 5408 10848 5424 10912
rect 5488 10848 5496 10912
rect 5176 10587 5496 10848
rect 5176 10351 5218 10587
rect 5454 10351 5496 10587
rect 5176 9824 5496 10351
rect 5176 9760 5184 9824
rect 5248 9760 5264 9824
rect 5328 9760 5344 9824
rect 5408 9760 5424 9824
rect 5488 9760 5496 9824
rect 5176 8736 5496 9760
rect 5176 8672 5184 8736
rect 5248 8672 5264 8736
rect 5328 8672 5344 8736
rect 5408 8672 5424 8736
rect 5488 8672 5496 8736
rect 5176 7648 5496 8672
rect 5176 7584 5184 7648
rect 5248 7584 5264 7648
rect 5328 7584 5344 7648
rect 5408 7584 5424 7648
rect 5488 7584 5496 7648
rect 5176 6560 5496 7584
rect 5176 6496 5184 6560
rect 5248 6496 5264 6560
rect 5328 6496 5344 6560
rect 5408 6496 5424 6560
rect 5488 6496 5496 6560
rect 5176 6416 5496 6496
rect 5176 6180 5218 6416
rect 5454 6180 5496 6416
rect 5176 5472 5496 6180
rect 5176 5408 5184 5472
rect 5248 5408 5264 5472
rect 5328 5408 5344 5472
rect 5408 5408 5424 5472
rect 5488 5408 5496 5472
rect 5176 4384 5496 5408
rect 5176 4320 5184 4384
rect 5248 4320 5264 4384
rect 5328 4320 5344 4384
rect 5408 4320 5424 4384
rect 5488 4320 5496 4384
rect 5176 3296 5496 4320
rect 5176 3232 5184 3296
rect 5248 3232 5264 3296
rect 5328 3232 5344 3296
rect 5408 3232 5424 3296
rect 5488 3232 5496 3296
rect 5176 2208 5496 3232
rect 5176 2144 5184 2208
rect 5248 2144 5264 2208
rect 5328 2144 5344 2208
rect 5408 2144 5424 2208
rect 5488 2144 5496 2208
rect 5176 2128 5496 2144
rect 7292 14720 7612 14736
rect 7292 14656 7300 14720
rect 7364 14656 7380 14720
rect 7444 14656 7460 14720
rect 7524 14656 7540 14720
rect 7604 14656 7612 14720
rect 7292 13632 7612 14656
rect 7292 13568 7300 13632
rect 7364 13568 7380 13632
rect 7444 13568 7460 13632
rect 7524 13568 7540 13632
rect 7604 13568 7612 13632
rect 7292 12672 7612 13568
rect 7292 12544 7334 12672
rect 7570 12544 7612 12672
rect 7292 12480 7300 12544
rect 7604 12480 7612 12544
rect 7292 12436 7334 12480
rect 7570 12436 7612 12480
rect 7292 11456 7612 12436
rect 7292 11392 7300 11456
rect 7364 11392 7380 11456
rect 7444 11392 7460 11456
rect 7524 11392 7540 11456
rect 7604 11392 7612 11456
rect 7292 10368 7612 11392
rect 7292 10304 7300 10368
rect 7364 10304 7380 10368
rect 7444 10304 7460 10368
rect 7524 10304 7540 10368
rect 7604 10304 7612 10368
rect 7292 9280 7612 10304
rect 7292 9216 7300 9280
rect 7364 9216 7380 9280
rect 7444 9216 7460 9280
rect 7524 9216 7540 9280
rect 7604 9216 7612 9280
rect 7292 8502 7612 9216
rect 7292 8266 7334 8502
rect 7570 8266 7612 8502
rect 7292 8192 7612 8266
rect 7292 8128 7300 8192
rect 7364 8128 7380 8192
rect 7444 8128 7460 8192
rect 7524 8128 7540 8192
rect 7604 8128 7612 8192
rect 7292 7104 7612 8128
rect 7292 7040 7300 7104
rect 7364 7040 7380 7104
rect 7444 7040 7460 7104
rect 7524 7040 7540 7104
rect 7604 7040 7612 7104
rect 7292 6016 7612 7040
rect 7292 5952 7300 6016
rect 7364 5952 7380 6016
rect 7444 5952 7460 6016
rect 7524 5952 7540 6016
rect 7604 5952 7612 6016
rect 7292 4928 7612 5952
rect 7292 4864 7300 4928
rect 7364 4864 7380 4928
rect 7444 4864 7460 4928
rect 7524 4864 7540 4928
rect 7604 4864 7612 4928
rect 7292 4331 7612 4864
rect 7292 4095 7334 4331
rect 7570 4095 7612 4331
rect 7292 3840 7612 4095
rect 7292 3776 7300 3840
rect 7364 3776 7380 3840
rect 7444 3776 7460 3840
rect 7524 3776 7540 3840
rect 7604 3776 7612 3840
rect 7292 2752 7612 3776
rect 7292 2688 7300 2752
rect 7364 2688 7380 2752
rect 7444 2688 7460 2752
rect 7524 2688 7540 2752
rect 7604 2688 7612 2752
rect 7292 2128 7612 2688
rect 9408 14176 9728 14736
rect 9408 14112 9416 14176
rect 9480 14112 9496 14176
rect 9560 14112 9576 14176
rect 9640 14112 9656 14176
rect 9720 14112 9728 14176
rect 9408 13088 9728 14112
rect 9408 13024 9416 13088
rect 9480 13024 9496 13088
rect 9560 13024 9576 13088
rect 9640 13024 9656 13088
rect 9720 13024 9728 13088
rect 9408 12000 9728 13024
rect 9408 11936 9416 12000
rect 9480 11936 9496 12000
rect 9560 11936 9576 12000
rect 9640 11936 9656 12000
rect 9720 11936 9728 12000
rect 9408 10912 9728 11936
rect 9408 10848 9416 10912
rect 9480 10848 9496 10912
rect 9560 10848 9576 10912
rect 9640 10848 9656 10912
rect 9720 10848 9728 10912
rect 9408 10587 9728 10848
rect 9408 10351 9450 10587
rect 9686 10351 9728 10587
rect 9408 9824 9728 10351
rect 9408 9760 9416 9824
rect 9480 9760 9496 9824
rect 9560 9760 9576 9824
rect 9640 9760 9656 9824
rect 9720 9760 9728 9824
rect 9408 8736 9728 9760
rect 9408 8672 9416 8736
rect 9480 8672 9496 8736
rect 9560 8672 9576 8736
rect 9640 8672 9656 8736
rect 9720 8672 9728 8736
rect 9408 7648 9728 8672
rect 9408 7584 9416 7648
rect 9480 7584 9496 7648
rect 9560 7584 9576 7648
rect 9640 7584 9656 7648
rect 9720 7584 9728 7648
rect 9408 6560 9728 7584
rect 9408 6496 9416 6560
rect 9480 6496 9496 6560
rect 9560 6496 9576 6560
rect 9640 6496 9656 6560
rect 9720 6496 9728 6560
rect 9408 6416 9728 6496
rect 9408 6180 9450 6416
rect 9686 6180 9728 6416
rect 9408 5472 9728 6180
rect 9408 5408 9416 5472
rect 9480 5408 9496 5472
rect 9560 5408 9576 5472
rect 9640 5408 9656 5472
rect 9720 5408 9728 5472
rect 9408 4384 9728 5408
rect 9408 4320 9416 4384
rect 9480 4320 9496 4384
rect 9560 4320 9576 4384
rect 9640 4320 9656 4384
rect 9720 4320 9728 4384
rect 9408 3296 9728 4320
rect 9408 3232 9416 3296
rect 9480 3232 9496 3296
rect 9560 3232 9576 3296
rect 9640 3232 9656 3296
rect 9720 3232 9728 3296
rect 9408 2208 9728 3232
rect 9408 2144 9416 2208
rect 9480 2144 9496 2208
rect 9560 2144 9576 2208
rect 9640 2144 9656 2208
rect 9720 2144 9728 2208
rect 9408 2128 9728 2144
rect 11524 14720 11844 14736
rect 11524 14656 11532 14720
rect 11596 14656 11612 14720
rect 11676 14656 11692 14720
rect 11756 14656 11772 14720
rect 11836 14656 11844 14720
rect 11524 13632 11844 14656
rect 11524 13568 11532 13632
rect 11596 13568 11612 13632
rect 11676 13568 11692 13632
rect 11756 13568 11772 13632
rect 11836 13568 11844 13632
rect 11524 12672 11844 13568
rect 11524 12544 11566 12672
rect 11802 12544 11844 12672
rect 11524 12480 11532 12544
rect 11836 12480 11844 12544
rect 11524 12436 11566 12480
rect 11802 12436 11844 12480
rect 11524 11456 11844 12436
rect 11524 11392 11532 11456
rect 11596 11392 11612 11456
rect 11676 11392 11692 11456
rect 11756 11392 11772 11456
rect 11836 11392 11844 11456
rect 11524 10368 11844 11392
rect 11524 10304 11532 10368
rect 11596 10304 11612 10368
rect 11676 10304 11692 10368
rect 11756 10304 11772 10368
rect 11836 10304 11844 10368
rect 11524 9280 11844 10304
rect 11524 9216 11532 9280
rect 11596 9216 11612 9280
rect 11676 9216 11692 9280
rect 11756 9216 11772 9280
rect 11836 9216 11844 9280
rect 11524 8502 11844 9216
rect 11524 8266 11566 8502
rect 11802 8266 11844 8502
rect 11524 8192 11844 8266
rect 11524 8128 11532 8192
rect 11596 8128 11612 8192
rect 11676 8128 11692 8192
rect 11756 8128 11772 8192
rect 11836 8128 11844 8192
rect 11524 7104 11844 8128
rect 11524 7040 11532 7104
rect 11596 7040 11612 7104
rect 11676 7040 11692 7104
rect 11756 7040 11772 7104
rect 11836 7040 11844 7104
rect 11524 6016 11844 7040
rect 11524 5952 11532 6016
rect 11596 5952 11612 6016
rect 11676 5952 11692 6016
rect 11756 5952 11772 6016
rect 11836 5952 11844 6016
rect 11524 4928 11844 5952
rect 11524 4864 11532 4928
rect 11596 4864 11612 4928
rect 11676 4864 11692 4928
rect 11756 4864 11772 4928
rect 11836 4864 11844 4928
rect 11524 4331 11844 4864
rect 11524 4095 11566 4331
rect 11802 4095 11844 4331
rect 11524 3840 11844 4095
rect 11524 3776 11532 3840
rect 11596 3776 11612 3840
rect 11676 3776 11692 3840
rect 11756 3776 11772 3840
rect 11836 3776 11844 3840
rect 11524 2752 11844 3776
rect 11524 2688 11532 2752
rect 11596 2688 11612 2752
rect 11676 2688 11692 2752
rect 11756 2688 11772 2752
rect 11836 2688 11844 2752
rect 11524 2128 11844 2688
<< via4 >>
rect 3102 12544 3338 12672
rect 3102 12480 3132 12544
rect 3132 12480 3148 12544
rect 3148 12480 3212 12544
rect 3212 12480 3228 12544
rect 3228 12480 3292 12544
rect 3292 12480 3308 12544
rect 3308 12480 3338 12544
rect 3102 12436 3338 12480
rect 3102 8266 3338 8502
rect 3102 4095 3338 4331
rect 5218 10351 5454 10587
rect 5218 6180 5454 6416
rect 7334 12544 7570 12672
rect 7334 12480 7364 12544
rect 7364 12480 7380 12544
rect 7380 12480 7444 12544
rect 7444 12480 7460 12544
rect 7460 12480 7524 12544
rect 7524 12480 7540 12544
rect 7540 12480 7570 12544
rect 7334 12436 7570 12480
rect 7334 8266 7570 8502
rect 7334 4095 7570 4331
rect 9450 10351 9686 10587
rect 9450 6180 9686 6416
rect 11566 12544 11802 12672
rect 11566 12480 11596 12544
rect 11596 12480 11612 12544
rect 11612 12480 11676 12544
rect 11676 12480 11692 12544
rect 11692 12480 11756 12544
rect 11756 12480 11772 12544
rect 11772 12480 11802 12544
rect 11566 12436 11802 12480
rect 11566 8266 11802 8502
rect 11566 4095 11802 4331
<< metal5 >>
rect 1104 12672 13800 12715
rect 1104 12436 3102 12672
rect 3338 12436 7334 12672
rect 7570 12436 11566 12672
rect 11802 12436 13800 12672
rect 1104 12394 13800 12436
rect 1104 10587 13800 10629
rect 1104 10351 5218 10587
rect 5454 10351 9450 10587
rect 9686 10351 13800 10587
rect 1104 10309 13800 10351
rect 1104 8502 13800 8544
rect 1104 8266 3102 8502
rect 3338 8266 7334 8502
rect 7570 8266 11566 8502
rect 11802 8266 13800 8502
rect 1104 8224 13800 8266
rect 1104 6416 13800 6459
rect 1104 6180 5218 6416
rect 5454 6180 9450 6416
rect 9686 6180 13800 6416
rect 1104 6138 13800 6180
rect 1104 4331 13800 4373
rect 1104 4095 3102 4331
rect 3338 4095 7334 4331
rect 7570 4095 11566 4331
rect 11802 4095 13800 4331
rect 1104 4053 13800 4095
use sky130_fd_sc_hd__decap_8  FILLER_0_7
timestamp 0
transform 1 0 1748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_61
timestamp 0
transform 1 0 6716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73
timestamp 0
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 0
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123
timestamp 0
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 0
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_7
timestamp 0
transform 1 0 1748 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 0
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_31
timestamp 0
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_43
timestamp 0
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 0
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 0
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_31
timestamp 0
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 0
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 0
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_37
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 0
transform 1 0 5152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 0
transform 1 0 6256 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 0
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 0
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 0
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_73
timestamp 0
transform 1 0 7820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_77
timestamp 0
transform 1 0 8188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_89
timestamp 0
transform 1 0 9292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_101
timestamp 0
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 0
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 0
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 0
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 0
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_36
timestamp 0
transform 1 0 4416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_59
timestamp 0
transform 1 0 6532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_88
timestamp 0
transform 1 0 9200 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_100
timestamp 0
transform 1 0 10304 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_112
timestamp 0
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_124
timestamp 0
transform 1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_132
timestamp 0
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_20
timestamp 0
transform 1 0 2944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 0
transform 1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 0
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 0
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_63
timestamp 0
transform 1 0 6900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 0
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_97
timestamp 0
transform 1 0 10028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 0
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp 0
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 0
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_36
timestamp 0
transform 1 0 4416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_45
timestamp 0
transform 1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 0
transform 1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_68
timestamp 0
transform 1 0 7360 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 0
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_101
timestamp 0
transform 1 0 10396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_113
timestamp 0
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_125
timestamp 0
transform 1 0 12604 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_13
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 0
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_31
timestamp 0
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp 0
transform 1 0 4968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 0
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_60
timestamp 0
transform 1 0 6624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_64
timestamp 0
transform 1 0 6992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 0
transform 1 0 8004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 0
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 0
transform 1 0 9752 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 0
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_131
timestamp 0
transform 1 0 13156 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 0
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_49
timestamp 0
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_69
timestamp 0
transform 1 0 7452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 0
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 0
transform 1 0 9660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 0
transform 1 0 10764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 0
transform 1 0 11868 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_129
timestamp 0
transform 1 0 12972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 0
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 0
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_43
timestamp 0
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 0
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_71
timestamp 0
transform 1 0 7636 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 0
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_87
timestamp 0
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_99
timestamp 0
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 0
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_10
timestamp 0
transform 1 0 2024 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 0
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_34
timestamp 0
transform 1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 0
transform 1 0 4968 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp 0
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_66
timestamp 0
transform 1 0 7176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_78
timestamp 0
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_89
timestamp 0
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_96
timestamp 0
transform 1 0 9936 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_108
timestamp 0
transform 1 0 11040 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_120
timestamp 0
transform 1 0 12144 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_132
timestamp 0
transform 1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_20
timestamp 0
transform 1 0 2944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 0
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_38
timestamp 0
transform 1 0 4600 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_44
timestamp 0
transform 1 0 5152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 0
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_64
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 0
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_85
timestamp 0
transform 1 0 8924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 0
transform 1 0 13340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 0
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_57
timestamp 0
transform 1 0 6348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 0
transform 1 0 6716 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_73
timestamp 0
transform 1 0 7820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 0
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_101
timestamp 0
transform 1 0 10396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_113
timestamp 0
transform 1 0 11500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_125
timestamp 0
transform 1 0 12604 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 0
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_44
timestamp 0
transform 1 0 5152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_48
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 0
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 0
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_74
timestamp 0
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 0
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 0
transform 1 0 10120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 0
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 0
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_6
timestamp 0
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 0
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 0
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_44
timestamp 0
transform 1 0 5152 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 0
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 0
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 0
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_65
timestamp 0
transform 1 0 7084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_77
timestamp 0
transform 1 0 8188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_89
timestamp 0
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 0
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 0
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 0
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 0
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp 0
transform 1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 0
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 0
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 0
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_131
timestamp 0
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_7
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 0
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_61
timestamp 0
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 0
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 0
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_91
timestamp 0
transform 1 0 9476 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_103
timestamp 0
transform 1 0 10580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 0
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_113
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_123
timestamp 0
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 0
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 13800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 13800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 13800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 13800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 13800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 13800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 13800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 13800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 13800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 13800 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 13800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 13800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 13800 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 13800 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 13800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 13800 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 0
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _063_
timestamp 0
transform 1 0 2392 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _064_
timestamp 0
transform -1 0 5060 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _065_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _066_
timestamp 0
transform -1 0 4968 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _067_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _068_
timestamp 0
transform 1 0 6900 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _069_
timestamp 0
transform -1 0 7912 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _070_
timestamp 0
transform -1 0 7084 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 0
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _072_
timestamp 0
transform -1 0 9108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 0
transform -1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _074_
timestamp 0
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _075_
timestamp 0
transform 1 0 1932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _076_
timestamp 0
transform 1 0 3312 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _077_
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _078_
timestamp 0
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 0
transform -1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _080_
timestamp 0
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _081_
timestamp 0
transform -1 0 3864 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _082_
timestamp 0
transform 1 0 2852 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _083_
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _084_
timestamp 0
transform -1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _085_
timestamp 0
transform -1 0 5244 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_
timestamp 0
transform -1 0 4600 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _087_
timestamp 0
transform -1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _088_
timestamp 0
transform 1 0 2668 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _089_
timestamp 0
transform 1 0 3036 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _090_
timestamp 0
transform -1 0 3312 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _091_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _092_
timestamp 0
transform -1 0 5336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _093_
timestamp 0
transform 1 0 4784 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _094_
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _095_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _096_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _097_
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _098_
timestamp 0
transform -1 0 8004 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _099_
timestamp 0
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _100_
timestamp 0
transform -1 0 5888 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _101_
timestamp 0
transform 1 0 9108 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _102_
timestamp 0
transform 1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _103_
timestamp 0
transform -1 0 6900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _104_
timestamp 0
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _105_
timestamp 0
transform 1 0 7728 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _106_
timestamp 0
transform 1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 0
transform 1 0 6256 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _108_
timestamp 0
transform 1 0 7360 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _109_
timestamp 0
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _110_
timestamp 0
transform 1 0 8372 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _111_
timestamp 0
transform 1 0 7820 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 0
transform 1 0 8280 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _115_
timestamp 0
transform -1 0 8372 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _116_
timestamp 0
transform -1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _117_
timestamp 0
transform -1 0 8280 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _118_
timestamp 0
transform -1 0 8464 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _119_
timestamp 0
transform 1 0 9568 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 0
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _121_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _122_
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _123_
timestamp 0
transform 1 0 6532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 0
transform 1 0 6440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _125_
timestamp 0
transform 1 0 5244 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _126_
timestamp 0
transform 1 0 4600 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  _127_
timestamp 0
transform 1 0 1748 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _128_
timestamp 0
transform -1 0 2944 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _129_
timestamp 0
transform 1 0 3680 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _130_
timestamp 0
transform 1 0 4140 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _131_
timestamp 0
transform 1 0 1472 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _132_
timestamp 0
transform -1 0 3956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _133_
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _134_
timestamp 0
transform 1 0 1472 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _135_
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _136_
timestamp 0
transform 1 0 6900 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _137_
timestamp 0
transform -1 0 10396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _138_
timestamp 0
transform -1 0 8740 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _139_
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _140_
timestamp 0
transform 1 0 9292 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _141_
timestamp 0
transform 1 0 5888 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _142_
timestamp 0
transform 1 0 4508 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 0
transform -1 0 13156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 0
transform -1 0 13156 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 0
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 0
transform -1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 0
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 0
transform 1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 0
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform 1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 3036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 0
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 0
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 0
transform -1 0 1748 0 1 14144
box -38 -48 406 592
<< labels >>
rlabel metal5 s 1104 6139 13800 6459 4 VGND
port 1 nsew
rlabel metal5 s 1104 10309 13800 10629 4 VGND
port 1 nsew
rlabel metal4 s 5176 2128 5496 14736 4 VGND
port 1 nsew
rlabel metal4 s 9408 2128 9728 14736 4 VGND
port 1 nsew
rlabel metal5 s 1104 4053 13800 4373 4 VPWR
port 2 nsew
rlabel metal5 s 1104 8224 13800 8544 4 VPWR
port 2 nsew
rlabel metal5 s 1104 12395 13800 12715 4 VPWR
port 2 nsew
rlabel metal4 s 3060 2128 3380 14736 4 VPWR
port 2 nsew
rlabel metal4 s 7292 2128 7612 14736 4 VPWR
port 2 nsew
rlabel metal4 s 11524 2128 11844 14736 4 VPWR
port 2 nsew
rlabel metal3 s 14181 3408 14981 3528 4 clock
port 3 nsew
rlabel metal2 s 14830 16325 14886 17125 4 count[0]
port 4 nsew
rlabel metal2 s 9034 16325 9090 17125 4 count[10]
port 5 nsew
rlabel metal2 s 5814 0 5870 800 4 count[11]
port 6 nsew
rlabel metal3 s 14181 13608 14981 13728 4 count[12]
port 7 nsew
rlabel metal3 s 14181 8 14981 128 4 count[13]
port 8 nsew
rlabel metal3 s 0 12928 800 13048 4 count[14]
port 9 nsew
rlabel metal2 s 5814 16325 5870 17125 4 count[15]
port 10 nsew
rlabel metal2 s 18 0 74 800 4 count[1]
port 11 nsew
rlabel metal2 s 2594 16325 2650 17125 4 count[2]
port 12 nsew
rlabel metal2 s 12254 0 12310 800 4 count[3]
port 13 nsew
rlabel metal2 s 2594 0 2650 800 4 count[4]
port 14 nsew
rlabel metal3 s 0 2728 800 2848 4 count[5]
port 15 nsew
rlabel metal3 s 14181 10208 14981 10328 4 count[6]
port 16 nsew
rlabel metal3 s 0 6128 800 6248 4 count[7]
port 17 nsew
rlabel metal2 s 12254 16325 12310 17125 4 count[8]
port 18 nsew
rlabel metal2 s 9034 0 9090 800 4 count[9]
port 19 nsew
rlabel metal3 s 0 9528 800 9648 4 count_en
port 20 nsew
rlabel metal3 s 0 16328 800 16448 4 count_tc
port 21 nsew
rlabel metal3 s 14181 6808 14981 6928 4 reset
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 14981 17125
<< end >>
